library verilog;
use verilog.vl_types.all;
entity flow is
    port(
        debug_valid     : out    vl_logic;
        debug_num_0     : out    vl_logic_vector(12 downto 0);
        debug_num_1     : out    vl_logic_vector(12 downto 0);
        debug_num_2     : out    vl_logic_vector(12 downto 0);
        debug_num_3     : out    vl_logic_vector(12 downto 0);
        debug_num_4     : out    vl_logic_vector(12 downto 0);
        debug_num_5     : out    vl_logic_vector(13 downto 0);
        debug_num_6     : out    vl_logic;
        debug_num_7     : out    vl_logic;
        debug_num_8     : out    vl_logic;
        t1              : in     vl_logic_vector(7 downto 0);
        t2              : in     vl_logic_vector(7 downto 0);
        t3              : in     vl_logic_vector(7 downto 0);
        b1              : in     vl_logic_vector(7 downto 0);
        b2              : in     vl_logic_vector(7 downto 0);
        b3              : in     vl_logic_vector(7 downto 0);
        i1              : in     vl_logic_vector(7 downto 0);
        i2              : in     vl_logic_vector(7 downto 0);
        i_clock         : in     vl_logic;
        i_reset         : in     vl_logic;
        i_valid         : in     vl_logic;
        i_mode          : in     vl_logic_vector(1 downto 0);
        i_row           : in     vl_logic_vector(7 downto 0);
        o_dir           : out    vl_logic_vector(2 downto 0);
        o_edge          : out    vl_logic;
        o_valid         : out    vl_logic;
        o_mode          : out    vl_logic_vector(1 downto 0);
        o_row           : out    vl_logic_vector(7 downto 0);
        p_ix258_ix248_nx13: out    vl_logic;
        p_ix258_ix249_nx13: out    vl_logic;
        p_ix258_ix250_nx13: out    vl_logic;
        p_ix258_ix251_nx13: out    vl_logic;
        p_ix258_ix252_nx13: out    vl_logic;
        p_ix258_ix253_nx13: out    vl_logic;
        p_ix258_ix254_nx13: out    vl_logic;
        p_ix258_ix255_nx13: out    vl_logic;
        p_not_rtlc5n47  : out    vl_logic;
        \p_p23_10_\     : out    vl_logic;
        \p_p23_9_\      : out    vl_logic;
        \p_p23_8_\      : out    vl_logic;
        \p_p23_7_\      : out    vl_logic;
        \p_p23_6_\      : out    vl_logic;
        \p_p23_5_\      : out    vl_logic;
        \p_p23_4_\      : out    vl_logic;
        \p_p23_3_\      : out    vl_logic;
        \p_p23_2_\      : out    vl_logic;
        \p_p23_1_\      : out    vl_logic;
        \p_p23_0_\      : out    vl_logic;
        \p_p21_4n0r2_12_\: out    vl_logic;
        \p_p21_4n0r2_11_\: out    vl_logic;
        \p_p21_4n0r2_10_\: out    vl_logic;
        \p_p21_4n0r2_9_\: out    vl_logic;
        \p_p21_4n0r2_8_\: out    vl_logic;
        \p_p21_4n0r2_7_\: out    vl_logic;
        \p_p21_4n0r2_6_\: out    vl_logic;
        \p_p21_4n0r2_5_\: out    vl_logic;
        \p_p21_4n0r2_4_\: out    vl_logic;
        \p_p21_4n0r2_3_\: out    vl_logic;
        \p_p21_4n0r2_2_\: out    vl_logic;
        \p_p21_4n0r2_1_\: out    vl_logic;
        \p_p21_4n0r3_0_\: out    vl_logic;
        \p_p22_4n0r2_12_\: out    vl_logic;
        \p_p22_4n0r2_11_\: out    vl_logic;
        \p_p22_4n0r2_10_\: out    vl_logic;
        \p_p22_4n0r2_9_\: out    vl_logic;
        \p_p22_4n0r2_8_\: out    vl_logic;
        \p_p22_4n0r2_7_\: out    vl_logic;
        \p_p22_4n0r2_6_\: out    vl_logic;
        \p_p22_4n0r2_5_\: out    vl_logic;
        \p_p22_4n0r2_4_\: out    vl_logic;
        \p_p22_4n0r2_3_\: out    vl_logic;
        \p_p22_4n0r2_2_\: out    vl_logic;
        \p_p22_4n0r2_1_\: out    vl_logic;
        \p_p22_4n0r3_0_\: out    vl_logic;
        \p_p5m_1_\      : out    vl_logic;
        \p_p5m_0_\      : out    vl_logic
    );
end flow;
