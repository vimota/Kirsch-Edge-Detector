
-- 
-- Definition of  kirsch
-- 
--      Sat Jul 19 23:39:09 2014
--      
--      Precision RTL Synthesis, 2008a.47
-- 

library IEEE;library altera_mf;library lpm;library altera; 
 use IEEE.STD_LOGIC_1164.ALL;
 use altera_mf.altera_mf_components.all, lpm.lpm_components.all, altera.altera_primitives_components.all;

entity ram_new_0_mem_8_8_main is 
   port (
      wr_data1 : IN std_logic_vector (7 DOWNTO 0) ;
      rd_data1 : OUT std_logic_vector (7 DOWNTO 0) ;
      addr1 : IN std_logic_vector (7 DOWNTO 0) ;
      wr_clk1 : IN std_logic ;
      rd_clk1 : IN std_logic ;
      wr_ena1 : IN std_logic ;
      rd_ena1 : IN std_logic ;
      ena1 : IN std_logic ;
      rst1 : IN std_logic ;
      regce1 : IN std_logic) ;
end ram_new_0_mem_8_8_main ;

architecture INTERFACE_unfold_2 of ram_new_0_mem_8_8_main is 
   procedure DFFPC (
      constant data   : in std_logic;
      constant preset : in std_logic;
      constant clear  : in std_logic;
      signal clk      : in std_logic;
      signal q        : out std_logic)
   is begin
       if (preset = '1') then
           q <= '1' ;
       elsif (clear = '1') then
           q <= '0' ;
       elsif (clk'event and clk'last_value = '0' and clk = '1') then
           q <= data and data ;    -- takes care of q<='X' if data='Z'
       end if ;
       if ((clear/='1' or preset/='1') and clk/='0' and clk/='1') then
           q <= 'X' ;
       end if ;
   end DFFPC ;
   component clocked_ram_8_8_256_F_T_F_F_F_F_F_F
      generic (ram_type : integer := 2;
         dual_addresses : string := "TRUE") ;
      
      port (
         clk : IN std_logic ;
         we : IN std_logic ;
         address : IN std_logic_vector (7 DOWNTO 0) ;
         data : IN std_logic_vector (7 DOWNTO 0) ;
         q : OUT std_logic_vector (7 DOWNTO 0) ;
         addr2 : IN std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   signal nx31, nx33, dup_0_reg_address_7, dup_0_reg_address_6, 
      dup_0_reg_address_5, dup_0_reg_address_4, dup_0_reg_address_3, 
      dup_0_reg_address_2, dup_0_reg_address_1, dup_0_reg_address_0, nx35, 
      nx37: std_logic ;

begin
   nx31 <= '0' ;
   nx33 <= '1' ;
   DFFPC (addr1(7),nx31,nx31,rd_clk1,dup_0_reg_address_7) ;
   DFFPC (addr1(6),nx31,nx31,rd_clk1,dup_0_reg_address_6) ;
   DFFPC (addr1(5),nx31,nx31,rd_clk1,dup_0_reg_address_5) ;
   DFFPC (addr1(4),nx31,nx31,rd_clk1,dup_0_reg_address_4) ;
   DFFPC (addr1(3),nx31,nx31,rd_clk1,dup_0_reg_address_3) ;
   DFFPC (addr1(2),nx31,nx31,rd_clk1,dup_0_reg_address_2) ;
   DFFPC (addr1(1),nx31,nx31,rd_clk1,dup_0_reg_address_1) ;
   DFFPC (addr1(0),nx31,nx31,rd_clk1,dup_0_reg_address_0) ;
   mem : clocked_ram_8_8_256_F_T_F_F_F_F_F_F port map ( clk=>wr_clk1, we=>
      nx35, address(7)=>addr1(7), address(6)=>addr1(6), address(5)=>addr1(5), 
      address(4)=>addr1(4), address(3)=>addr1(3), address(2)=>addr1(2), 
      address(1)=>addr1(1), address(0)=>addr1(0), data(7)=>wr_data1(7), 
      data(6)=>wr_data1(6), data(5)=>wr_data1(5), data(4)=>wr_data1(4), 
      data(3)=>wr_data1(3), data(2)=>wr_data1(2), data(1)=>wr_data1(1), 
      data(0)=>wr_data1(0), q(7)=>rd_data1(7), q(6)=>rd_data1(6), q(5)=>
      rd_data1(5), q(4)=>rd_data1(4), q(3)=>rd_data1(3), q(2)=>rd_data1(2), 
      q(1)=>rd_data1(1), q(0)=>rd_data1(0), addr2(7)=>dup_0_reg_address_7, 
      addr2(6)=>dup_0_reg_address_6, addr2(5)=>dup_0_reg_address_5, addr2(4)
      =>dup_0_reg_address_4, addr2(3)=>dup_0_reg_address_3, addr2(2)=>
      dup_0_reg_address_2, addr2(1)=>dup_0_reg_address_1, addr2(0)=>
      dup_0_reg_address_0);
   nx35 <= wr_ena1 AND ena1 ;
   nx37 <= rd_ena1 AND ena1 ;
end INTERFACE_unfold_2 ;

library IEEE;library altera_mf;library lpm;library altera; 
 use IEEE.STD_LOGIC_1164.ALL;
 use altera_mf.altera_mf_components.all, lpm.lpm_components.all, altera.altera_primitives_components.all;

entity mem_8_8 is 
   port (
      address : IN std_logic_vector (7 DOWNTO 0) ;
      clock : IN std_logic ;
      data : IN std_logic_vector (7 DOWNTO 0) ;
      wren : IN std_logic ;
      q : OUT std_logic_vector (7 DOWNTO 0)) ;
end mem_8_8 ;

architecture main_unfold_1 of mem_8_8 is 
   component ram_new_0_mem_8_8_main
      port (
         wr_data1 : IN std_logic_vector (7 DOWNTO 0) ;
         rd_data1 : OUT std_logic_vector (7 DOWNTO 0) ;
         addr1 : IN std_logic_vector (7 DOWNTO 0) ;
         wr_clk1 : IN std_logic ;
         rd_clk1 : IN std_logic ;
         wr_ena1 : IN std_logic ;
         rd_ena1 : IN std_logic ;
         ena1 : IN std_logic ;
         rst1 : IN std_logic ;
         regce1 : IN std_logic) ;
   end component ;
   for mem : ram_new_0_mem_8_8_main use entity work.ram_new_0_mem_8_8_main(
   INTERFACE_unfold_2);
   signal GND, nx25: std_logic ;

begin
   GND <= '0' ;
   mem : ram_new_0_mem_8_8_main port map ( wr_data1(7)=>data(7), wr_data1(6)
      =>data(6), wr_data1(5)=>data(5), wr_data1(4)=>data(4), wr_data1(3)=>
      data(3), wr_data1(2)=>data(2), wr_data1(1)=>data(1), wr_data1(0)=>
      data(0), rd_data1(7)=>q(7), rd_data1(6)=>q(6), rd_data1(5)=>q(5), 
      rd_data1(4)=>q(4), rd_data1(3)=>q(3), rd_data1(2)=>q(2), rd_data1(1)=>
      q(1), rd_data1(0)=>q(0), addr1(7)=>address(7), addr1(6)=>address(6), 
      addr1(5)=>address(5), addr1(4)=>address(4), addr1(3)=>address(3), 
      addr1(2)=>address(2), addr1(1)=>address(1), addr1(0)=>address(0), 
      wr_clk1=>clock, rd_clk1=>clock, wr_ena1=>wren, rd_ena1=>nx25, ena1=>
      nx25, rst1=>GND, regce1=>nx25);
   nx25 <= '1' ;
end main_unfold_1 ;


architecture INTERFACE of ram_new_0_mem_8_8_main is 
   procedure DFFPC (
      constant data   : in std_logic;
      constant preset : in std_logic;
      constant clear  : in std_logic;
      signal clk      : in std_logic;
      signal q        : out std_logic)
   is begin
       if (preset = '1') then
           q <= '1' ;
       elsif (clear = '1') then
           q <= '0' ;
       elsif (clk'event and clk'last_value = '0' and clk = '1') then
           q <= data and data ;    -- takes care of q<='X' if data='Z'
       end if ;
       if ((clear/='1' or preset/='1') and clk/='0' and clk/='1') then
           q <= 'X' ;
       end if ;
   end DFFPC ;
   component clocked_ram_8_8_256_F_T_F_F_F_F_F_F
      generic (ram_type : integer := 2;
         dual_addresses : string := "TRUE") ;
      
      port (
         clk : IN std_logic ;
         we : IN std_logic ;
         address : IN std_logic_vector (7 DOWNTO 0) ;
         data : IN std_logic_vector (7 DOWNTO 0) ;
         q : OUT std_logic_vector (7 DOWNTO 0) ;
         addr2 : IN std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   signal nx31, nx33, dup_0_reg_address_7, dup_0_reg_address_6, 
      dup_0_reg_address_5, dup_0_reg_address_4, dup_0_reg_address_3, 
      dup_0_reg_address_2, dup_0_reg_address_1, dup_0_reg_address_0, nx35, 
      nx37: std_logic ;

begin
   nx31 <= '0' ;
   nx33 <= '1' ;
   DFFPC (addr1(7),nx31,nx31,rd_clk1,dup_0_reg_address_7) ;
   DFFPC (addr1(6),nx31,nx31,rd_clk1,dup_0_reg_address_6) ;
   DFFPC (addr1(5),nx31,nx31,rd_clk1,dup_0_reg_address_5) ;
   DFFPC (addr1(4),nx31,nx31,rd_clk1,dup_0_reg_address_4) ;
   DFFPC (addr1(3),nx31,nx31,rd_clk1,dup_0_reg_address_3) ;
   DFFPC (addr1(2),nx31,nx31,rd_clk1,dup_0_reg_address_2) ;
   DFFPC (addr1(1),nx31,nx31,rd_clk1,dup_0_reg_address_1) ;
   DFFPC (addr1(0),nx31,nx31,rd_clk1,dup_0_reg_address_0) ;
   mem : clocked_ram_8_8_256_F_T_F_F_F_F_F_F port map ( clk=>wr_clk1, we=>
      nx35, address(7)=>addr1(7), address(6)=>addr1(6), address(5)=>addr1(5), 
      address(4)=>addr1(4), address(3)=>addr1(3), address(2)=>addr1(2), 
      address(1)=>addr1(1), address(0)=>addr1(0), data(7)=>wr_data1(7), 
      data(6)=>wr_data1(6), data(5)=>wr_data1(5), data(4)=>wr_data1(4), 
      data(3)=>wr_data1(3), data(2)=>wr_data1(2), data(1)=>wr_data1(1), 
      data(0)=>wr_data1(0), q(7)=>rd_data1(7), q(6)=>rd_data1(6), q(5)=>
      rd_data1(5), q(4)=>rd_data1(4), q(3)=>rd_data1(3), q(2)=>rd_data1(2), 
      q(1)=>rd_data1(1), q(0)=>rd_data1(0), addr2(7)=>dup_0_reg_address_7, 
      addr2(6)=>dup_0_reg_address_6, addr2(5)=>dup_0_reg_address_5, addr2(4)
      =>dup_0_reg_address_4, addr2(3)=>dup_0_reg_address_3, addr2(2)=>
      dup_0_reg_address_2, addr2(1)=>dup_0_reg_address_1, addr2(0)=>
      dup_0_reg_address_0);
   nx35 <= wr_ena1 AND ena1 ;
   nx37 <= rd_ena1 AND ena1 ;
end INTERFACE ;


architecture main_unfold_2 of mem_8_8 is 
   component ram_new_0_mem_8_8_main
      port (
         wr_data1 : IN std_logic_vector (7 DOWNTO 0) ;
         rd_data1 : OUT std_logic_vector (7 DOWNTO 0) ;
         addr1 : IN std_logic_vector (7 DOWNTO 0) ;
         wr_clk1 : IN std_logic ;
         rd_clk1 : IN std_logic ;
         wr_ena1 : IN std_logic ;
         rd_ena1 : IN std_logic ;
         ena1 : IN std_logic ;
         rst1 : IN std_logic ;
         regce1 : IN std_logic) ;
   end component ;
   for mem : ram_new_0_mem_8_8_main use entity work.ram_new_0_mem_8_8_main(
   INTERFACE);
   signal GND, nx25: std_logic ;

begin
   GND <= '0' ;
   mem : ram_new_0_mem_8_8_main port map ( wr_data1(7)=>data(7), wr_data1(6)
      =>data(6), wr_data1(5)=>data(5), wr_data1(4)=>data(4), wr_data1(3)=>
      data(3), wr_data1(2)=>data(2), wr_data1(1)=>data(1), wr_data1(0)=>
      data(0), rd_data1(7)=>q(7), rd_data1(6)=>q(6), rd_data1(5)=>q(5), 
      rd_data1(4)=>q(4), rd_data1(3)=>q(3), rd_data1(2)=>q(2), rd_data1(1)=>
      q(1), rd_data1(0)=>q(0), addr1(7)=>address(7), addr1(6)=>address(6), 
      addr1(5)=>address(5), addr1(4)=>address(4), addr1(3)=>address(3), 
      addr1(2)=>address(2), addr1(1)=>address(1), addr1(0)=>address(0), 
      wr_clk1=>clock, rd_clk1=>clock, wr_ena1=>wren, rd_ena1=>nx25, ena1=>
      nx25, rst1=>GND, regce1=>nx25);
   nx25 <= '1' ;
end main_unfold_2 ;


architecture INTERFACE_unfold_1 of ram_new_0_mem_8_8_main is 
   procedure DFFPC (
      constant data   : in std_logic;
      constant preset : in std_logic;
      constant clear  : in std_logic;
      signal clk      : in std_logic;
      signal q        : out std_logic)
   is begin
       if (preset = '1') then
           q <= '1' ;
       elsif (clear = '1') then
           q <= '0' ;
       elsif (clk'event and clk'last_value = '0' and clk = '1') then
           q <= data and data ;    -- takes care of q<='X' if data='Z'
       end if ;
       if ((clear/='1' or preset/='1') and clk/='0' and clk/='1') then
           q <= 'X' ;
       end if ;
   end DFFPC ;
   component clocked_ram_8_8_256_F_T_F_F_F_F_F_F
      generic (ram_type : integer := 2;
         dual_addresses : string := "TRUE") ;
      
      port (
         clk : IN std_logic ;
         we : IN std_logic ;
         address : IN std_logic_vector (7 DOWNTO 0) ;
         data : IN std_logic_vector (7 DOWNTO 0) ;
         q : OUT std_logic_vector (7 DOWNTO 0) ;
         addr2 : IN std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   signal nx31, nx33, dup_0_reg_address_7, dup_0_reg_address_6, 
      dup_0_reg_address_5, dup_0_reg_address_4, dup_0_reg_address_3, 
      dup_0_reg_address_2, dup_0_reg_address_1, dup_0_reg_address_0, nx35, 
      nx37: std_logic ;

begin
   nx31 <= '0' ;
   nx33 <= '1' ;
   DFFPC (addr1(7),nx31,nx31,rd_clk1,dup_0_reg_address_7) ;
   DFFPC (addr1(6),nx31,nx31,rd_clk1,dup_0_reg_address_6) ;
   DFFPC (addr1(5),nx31,nx31,rd_clk1,dup_0_reg_address_5) ;
   DFFPC (addr1(4),nx31,nx31,rd_clk1,dup_0_reg_address_4) ;
   DFFPC (addr1(3),nx31,nx31,rd_clk1,dup_0_reg_address_3) ;
   DFFPC (addr1(2),nx31,nx31,rd_clk1,dup_0_reg_address_2) ;
   DFFPC (addr1(1),nx31,nx31,rd_clk1,dup_0_reg_address_1) ;
   DFFPC (addr1(0),nx31,nx31,rd_clk1,dup_0_reg_address_0) ;
   mem : clocked_ram_8_8_256_F_T_F_F_F_F_F_F port map ( clk=>wr_clk1, we=>
      nx35, address(7)=>addr1(7), address(6)=>addr1(6), address(5)=>addr1(5), 
      address(4)=>addr1(4), address(3)=>addr1(3), address(2)=>addr1(2), 
      address(1)=>addr1(1), address(0)=>addr1(0), data(7)=>wr_data1(7), 
      data(6)=>wr_data1(6), data(5)=>wr_data1(5), data(4)=>wr_data1(4), 
      data(3)=>wr_data1(3), data(2)=>wr_data1(2), data(1)=>wr_data1(1), 
      data(0)=>wr_data1(0), q(7)=>rd_data1(7), q(6)=>rd_data1(6), q(5)=>
      rd_data1(5), q(4)=>rd_data1(4), q(3)=>rd_data1(3), q(2)=>rd_data1(2), 
      q(1)=>rd_data1(1), q(0)=>rd_data1(0), addr2(7)=>dup_0_reg_address_7, 
      addr2(6)=>dup_0_reg_address_6, addr2(5)=>dup_0_reg_address_5, addr2(4)
      =>dup_0_reg_address_4, addr2(3)=>dup_0_reg_address_3, addr2(2)=>
      dup_0_reg_address_2, addr2(1)=>dup_0_reg_address_1, addr2(0)=>
      dup_0_reg_address_0);
   nx35 <= wr_ena1 AND ena1 ;
   nx37 <= rd_ena1 AND ena1 ;
end INTERFACE_unfold_1 ;


architecture main of mem_8_8 is 
   component ram_new_0_mem_8_8_main
      port (
         wr_data1 : IN std_logic_vector (7 DOWNTO 0) ;
         rd_data1 : OUT std_logic_vector (7 DOWNTO 0) ;
         addr1 : IN std_logic_vector (7 DOWNTO 0) ;
         wr_clk1 : IN std_logic ;
         rd_clk1 : IN std_logic ;
         wr_ena1 : IN std_logic ;
         rd_ena1 : IN std_logic ;
         ena1 : IN std_logic ;
         rst1 : IN std_logic ;
         regce1 : IN std_logic) ;
   end component ;
   for mem : ram_new_0_mem_8_8_main use entity work.ram_new_0_mem_8_8_main(
   INTERFACE_unfold_1);
   signal GND, nx25: std_logic ;

begin
   GND <= '0' ;
   mem : ram_new_0_mem_8_8_main port map ( wr_data1(7)=>data(7), wr_data1(6)
      =>data(6), wr_data1(5)=>data(5), wr_data1(4)=>data(4), wr_data1(3)=>
      data(3), wr_data1(2)=>data(2), wr_data1(1)=>data(1), wr_data1(0)=>
      data(0), rd_data1(7)=>q(7), rd_data1(6)=>q(6), rd_data1(5)=>q(5), 
      rd_data1(4)=>q(4), rd_data1(3)=>q(3), rd_data1(2)=>q(2), rd_data1(1)=>
      q(1), rd_data1(0)=>q(0), addr1(7)=>address(7), addr1(6)=>address(6), 
      addr1(5)=>address(5), addr1(4)=>address(4), addr1(3)=>address(3), 
      addr1(2)=>address(2), addr1(1)=>address(1), addr1(0)=>address(0), 
      wr_clk1=>clock, rd_clk1=>clock, wr_ena1=>wren, rd_ena1=>nx25, ena1=>
      nx25, rst1=>GND, regce1=>nx25);
   nx25 <= '1' ;
end main ;

library IEEE;library altera_mf;library lpm;library altera; 
 use IEEE.STD_LOGIC_1164.ALL;
 use altera_mf.altera_mf_components.all, lpm.lpm_components.all, altera.altera_primitives_components.all;

entity counter_up_cnt_en_clock_0_8 is 
   port (
      clock : IN std_logic ;
      q : OUT std_logic_vector (7 DOWNTO 0) ;
      clk_en : IN std_logic ;
      aclear : IN std_logic ;
      sload : IN std_logic ;
      data : IN std_logic_vector (7 DOWNTO 0) ;
      aset : IN std_logic ;
      sclear : IN std_logic ;
      updn : IN std_logic ;
      cnt_en : IN std_logic) ;
end counter_up_cnt_en_clock_0_8 ;

architecture INTERFACE of counter_up_cnt_en_clock_0_8 is 
   procedure DFFPCE (
      constant data   : in std_logic;
      constant preset : in std_logic;
      constant clear  : in std_logic;
      constant enable : in std_logic;
      signal clk      : in std_logic;
      signal q        : out std_logic)
   is begin
       if (preset = '1') then
           q <= '1' ;
       elsif (clear = '1') then
           q <= '0' ;
       elsif (clk'event and clk'last_value = '0' and clk = '1') then
           if (enable = '1') then
               q <= data and data ;    -- takes care of q<='X' if data='Z'
           end if ;
       end if ;
       if ((clear/='1' or preset/='1') and clk/='0' and clk/='1') then
           q <= 'X' ;
       end if ;
   end DFFPCE ;
   component inc_8u_8u_0_0
      port (
         cin : IN std_logic ;
         a : IN std_logic_vector (7 DOWNTO 0) ;
         d : OUT std_logic_vector (7 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal GND, nx20, nx21, nx22, nx23, nx24, nx25, nx26, nx27, nx28, nx29, 
      nx30, nx31, nx32, nx33, nx34, nx35, PWR: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   q(7) <= nx21 ;
   q(6) <= nx23 ;
   q(5) <= nx25 ;
   q(4) <= nx27 ;
   q(3) <= nx29 ;
   q(2) <= nx31 ;
   q(1) <= nx33 ;
   q(0) <= nx35 ;
   GND <= '0' ;
   DFFPCE (nx20,GND,GND,cnt_en,clock,nx21) ;
   DFFPCE (nx22,GND,GND,cnt_en,clock,nx23) ;
   DFFPCE (nx24,GND,GND,cnt_en,clock,nx25) ;
   DFFPCE (nx26,GND,GND,cnt_en,clock,nx27) ;
   DFFPCE (nx28,GND,GND,cnt_en,clock,nx29) ;
   DFFPCE (nx30,GND,GND,cnt_en,clock,nx31) ;
   DFFPCE (nx32,GND,GND,cnt_en,clock,nx33) ;
   DFFPCE (nx34,GND,GND,cnt_en,clock,nx35) ;
   inc : inc_8u_8u_0_0 port map ( cin=>PWR, a(7)=>nx21, a(6)=>nx23, a(5)=>
      nx25, a(4)=>nx27, a(3)=>nx29, a(2)=>nx31, a(1)=>nx33, a(0)=>nx35, d(7)
      =>nx20, d(6)=>nx22, d(5)=>nx24, d(4)=>nx26, d(3)=>nx28, d(2)=>nx30, 
      d(1)=>nx32, d(0)=>nx34, cout=>DANGLING(0));
   PWR <= '1' ;
end INTERFACE ;

library IEEE;library altera_mf;library lpm;library altera; 
 use IEEE.STD_LOGIC_1164.ALL;
 use altera_mf.altera_mf_components.all, lpm.lpm_components.all, altera.altera_primitives_components.all;

entity counter_up_sclear_clock_clk_en_0_8 is 
   port (
      clock : IN std_logic ;
      q : OUT std_logic_vector (7 DOWNTO 0) ;
      clk_en : IN std_logic ;
      aclear : IN std_logic ;
      sload : IN std_logic ;
      data : IN std_logic_vector (7 DOWNTO 0) ;
      aset : IN std_logic ;
      sclear : IN std_logic ;
      updn : IN std_logic ;
      cnt_en : IN std_logic) ;
end counter_up_sclear_clock_clk_en_0_8 ;

architecture INTERFACE of counter_up_sclear_clock_clk_en_0_8 is 
   procedure DFFPCE (
      constant data   : in std_logic;
      constant preset : in std_logic;
      constant clear  : in std_logic;
      constant enable : in std_logic;
      signal clk      : in std_logic;
      signal q        : out std_logic)
   is begin
       if (preset = '1') then
           q <= '1' ;
       elsif (clear = '1') then
           q <= '0' ;
       elsif (clk'event and clk'last_value = '0' and clk = '1') then
           if (enable = '1') then
               q <= data and data ;    -- takes care of q<='X' if data='Z'
           end if ;
       end if ;
       if ((clear/='1' or preset/='1') and clk/='0' and clk/='1') then
           q <= 'X' ;
       end if ;
   end DFFPCE ;
   component inc_8u_8u_0_0
      port (
         cin : IN std_logic ;
         a : IN std_logic_vector (7 DOWNTO 0) ;
         d : OUT std_logic_vector (7 DOWNTO 0) ;
         cout : OUT std_logic) ;
   end component ;
   signal GND, nx20, nx21, nx22, nx23, nx24, nx25, nx26, nx27, nx28, nx29, 
      nx30, nx31, nx32, nx33, nx34, nx35, nx36, nx37, nx38, nx39, nx40, nx41, 
      nx42, nx43, PWR, NOT_SCLEAR: std_logic ;
   
   signal DANGLING : std_logic_vector (0 downto 0 );

begin
   q(7) <= nx21 ;
   q(6) <= nx23 ;
   q(5) <= nx25 ;
   q(4) <= nx27 ;
   q(3) <= nx29 ;
   q(2) <= nx31 ;
   q(1) <= nx33 ;
   q(0) <= nx35 ;
   GND <= '0' ;
   DFFPCE (nx20,GND,GND,clk_en,clock,nx21) ;
   DFFPCE (nx22,GND,GND,clk_en,clock,nx23) ;
   DFFPCE (nx24,GND,GND,clk_en,clock,nx25) ;
   DFFPCE (nx26,GND,GND,clk_en,clock,nx27) ;
   DFFPCE (nx28,GND,GND,clk_en,clock,nx29) ;
   DFFPCE (nx30,GND,GND,clk_en,clock,nx31) ;
   DFFPCE (nx32,GND,GND,clk_en,clock,nx33) ;
   DFFPCE (nx34,GND,GND,clk_en,clock,nx35) ;
   inc : inc_8u_8u_0_0 port map ( cin=>PWR, a(7)=>nx21, a(6)=>nx23, a(5)=>
      nx25, a(4)=>nx27, a(3)=>nx29, a(2)=>nx31, a(1)=>nx33, a(0)=>nx35, d(7)
      =>nx36, d(6)=>nx37, d(5)=>nx38, d(4)=>nx39, d(3)=>nx40, d(2)=>nx41, 
      d(1)=>nx42, d(0)=>nx43, cout=>DANGLING(0));
   PWR <= '1' ;
   NOT_SCLEAR <= NOT sclear ;
   nx20 <= nx36 AND NOT_SCLEAR ;
   nx22 <= nx37 AND NOT_SCLEAR ;
   nx24 <= nx38 AND NOT_SCLEAR ;
   nx26 <= nx39 AND NOT_SCLEAR ;
   nx28 <= nx40 AND NOT_SCLEAR ;
   nx30 <= nx41 AND NOT_SCLEAR ;
   nx32 <= nx42 AND NOT_SCLEAR ;
   nx34 <= nx43 AND NOT_SCLEAR ;
end INTERFACE ;

library IEEE;library altera_mf;library lpm;library altera; 
 use IEEE.STD_LOGIC_1164.ALL;
 use altera_mf.altera_mf_components.all, lpm.lpm_components.all, altera.altera_primitives_components.all;

entity memory_notri is 
   port (
      p_o_image0_9_7 : OUT std_logic_vector (1 DOWNTO 0) ;
      p_o_image0_9_1 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image0_9_2 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image0_9_3 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image0_9_4 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image0_9_5 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image0_9_6 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image0_8_7 : OUT std_logic_vector (1 DOWNTO 0) ;
      p_o_image0_8_1 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image0_8_2 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image0_8_3 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image0_8_4 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image0_8_5 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image0_8_6 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image0_7 : OUT std_logic_vector (2 DOWNTO 1) ;
      p_o_image0_1 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image0_2 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image0_3 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image0_4 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image0_5 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image0_6 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image1_9_7 : OUT std_logic_vector (1 DOWNTO 0) ;
      p_o_image1_9_1 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image1_9_2 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image1_9_3 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image1_9_4 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image1_9_5 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image1_9_6 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image1_8_7 : OUT std_logic_vector (1 DOWNTO 0) ;
      p_o_image1_8_1 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image1_8_2 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image1_8_3 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image1_8_4 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image1_8_5 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image1_8_6 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image1_7 : OUT std_logic_vector (2 DOWNTO 1) ;
      p_o_image1_1 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image1_2 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image1_3 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image1_4 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image1_5 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image1_6 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image2_9_7 : OUT std_logic_vector (1 DOWNTO 0) ;
      p_o_image2_9_1 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image2_9_2 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image2_9_3 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image2_9_4 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image2_9_5 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image2_9_6 : OUT std_logic_vector (0 DOWNTO 0) ;
      p_o_image2_8_7 : OUT std_logic_vector (1 DOWNTO 0) ;
      p_o_image2_8_1 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image2_8_2 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image2_8_3 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image2_8_4 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image2_8_5 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image2_8_6 : OUT std_logic_vector (1 DOWNTO 1) ;
      p_o_image2_7 : OUT std_logic_vector (2 DOWNTO 1) ;
      p_o_image2_1 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image2_2 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image2_3 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image2_4 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image2_5 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_o_image2_6 : OUT std_logic_vector (2 DOWNTO 2) ;
      p_i_pixel : IN std_logic_vector (7 DOWNTO 0) ;
      p_o_row : OUT std_logic_vector (7 DOWNTO 0) ;
      p_i_valid_rtlc_32_or_1 : IN std_logic_vector (2 DOWNTO 2) ;
      p_i_clock : IN std_logic ;
      p_o_column : OUT std_logic_vector (7 DOWNTO 0)) ;
end memory_notri ;

architecture main_unfold_1492 of memory_notri is 
   component mem_8_8
      port (
         address : IN std_logic_vector (7 DOWNTO 0) ;
         clock : IN std_logic ;
         data : IN std_logic_vector (7 DOWNTO 0) ;
         wren : IN std_logic ;
         q : OUT std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   component or_7u_7u
      port (
         a : IN std_logic_vector (6 DOWNTO 0) ;
         d : OUT std_logic) ;
   end component ;
   component or_3u_3u
      port (
         a : IN std_logic_vector (2 DOWNTO 0) ;
         d : OUT std_logic) ;
   end component ;
   component select_3_3
      port (
         a : IN std_logic_vector (2 DOWNTO 0) ;
         b : IN std_logic_vector (2 DOWNTO 0) ;
         d : OUT std_logic) ;
   end component ;
   component and_8u_8u
      port (
         a : IN std_logic_vector (7 DOWNTO 0) ;
         d : OUT std_logic) ;
   end component ;
   component counter_up_cnt_en_clock_0_8
      port (
         clock : IN std_logic ;
         q : OUT std_logic_vector (7 DOWNTO 0) ;
         clk_en : IN std_logic ;
         aclear : IN std_logic ;
         sload : IN std_logic ;
         data : IN std_logic_vector (7 DOWNTO 0) ;
         aset : IN std_logic ;
         sclear : IN std_logic ;
         updn : IN std_logic ;
         cnt_en : IN std_logic) ;
   end component ;
   component counter_up_sclear_clock_clk_en_0_8
      port (
         clock : IN std_logic ;
         q : OUT std_logic_vector (7 DOWNTO 0) ;
         clk_en : IN std_logic ;
         aclear : IN std_logic ;
         sload : IN std_logic ;
         data : IN std_logic_vector (7 DOWNTO 0) ;
         aset : IN std_logic ;
         sclear : IN std_logic ;
         updn : IN std_logic ;
         cnt_en : IN std_logic) ;
   end component ;
   procedure DFFPCE (
      constant data   : in std_logic;
      constant preset : in std_logic;
      constant clear  : in std_logic;
      constant enable : in std_logic;
      signal clk      : in std_logic;
      signal q        : out std_logic)
   is begin
       if (preset = '1') then
           q <= '1' ;
       elsif (clear = '1') then
           q <= '0' ;
       elsif (clk'event and clk'last_value = '0' and clk = '1') then
           if (enable = '1') then
               q <= data and data ;    -- takes care of q<='X' if data='Z'
           end if ;
       end if ;
       if ((clear/='1' or preset/='1') and clk/='0' and clk/='1') then
           q <= 'X' ;
       end if ;
   end DFFPCE ;
   procedure DFFPC (
      constant data   : in std_logic;
      constant preset : in std_logic;
      constant clear  : in std_logic;
      signal clk      : in std_logic;
      signal q        : out std_logic)
   is begin
       if (preset = '1') then
           q <= '1' ;
       elsif (clear = '1') then
           q <= '0' ;
       elsif (clk'event and clk'last_value = '0' and clk = '1') then
           q <= data and data ;    -- takes care of q<='X' if data='Z'
       end if ;
       if ((clear/='1' or preset/='1') and clk/='0' and clk/='1') then
           q <= 'X' ;
       end if ;
   end DFFPC ;
   for u_mem1 : mem_8_8 use entity work.mem_8_8(main_unfold_1);
   for u_mem2 : mem_8_8 use entity work.mem_8_8(main_unfold_2);
   for u_mem3 : mem_8_8 use entity work.mem_8_8(main);
   signal o_image1_0_7_rename21: std_logic_vector (1 DOWNTO 0) ;
   
   signal o_image1_0_1_rename22: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image1_0_2_rename23: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image1_0_3_rename24: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image1_0_4_rename25: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image1_0_5_rename26: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image1_0_6_rename27: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image1_1_7_rename28: std_logic_vector (1 DOWNTO 0) ;
   
   signal o_image1_1_1_rename29: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image1_1_2_rename30: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image1_1_3_rename31: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image1_1_4_rename32: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image1_1_5_rename33: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image1_1_6_rename34: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image1_2_7_rename35: std_logic_vector (2 DOWNTO 1) ;
   
   signal o_image1_2_1_rename36: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image1_2_2_rename37: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image1_2_3_rename38: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image1_2_4_rename39: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image1_2_5_rename40: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image1_2_6_rename41: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image2_0_7_rename42: std_logic_vector (1 DOWNTO 0) ;
   
   signal o_image2_0_1_rename43: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image2_0_2_rename44: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image2_0_3_rename45: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image2_0_4_rename46: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image2_0_5_rename47: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image2_0_6_rename48: std_logic_vector (0 DOWNTO 0) ;
   
   signal o_image2_1_7_rename49: std_logic_vector (1 DOWNTO 0) ;
   
   signal o_image2_1_1_rename50: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image2_1_2_rename51: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image2_1_3_rename52: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image2_1_4_rename53: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image2_1_5_rename54: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image2_1_6_rename55: std_logic_vector (1 DOWNTO 1) ;
   
   signal o_image2_2_7_rename56: std_logic_vector (2 DOWNTO 1) ;
   
   signal o_image2_2_1_rename57: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image2_2_2_rename58: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image2_2_3_rename59: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image2_2_4_rename60: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image2_2_5_rename61: std_logic_vector (2 DOWNTO 2) ;
   
   signal o_image2_2_6_rename62: std_logic_vector (2 DOWNTO 2) ;
   
   signal rtlcn234, rtlcn233, rtlcn231, rtlcn229, not_rtlc0n225: std_logic
    ;
   
   signal mem_wrn_current_0n4ss1: std_logic_vector (2 DOWNTO 0) ;
   
   signal first_bubble, not_rtlc0n172: std_logic ;
   
   signal buffer2_1n3ss1: std_logic_vector (23 DOWNTO 0) ;
   
   signal rtlc0n172, rtlcn226, rtlcn225, rtlcn217, rtlcn121, not_rtlcn226: 
   std_logic ;
   
   signal buffer2_1n1ss1: std_logic_vector (7 DOWNTO 0) ;
   
   signal rtlcn97, not_rtlcn225, rtlc1n272, o_row_7, o_row_6, o_row_5, 
      o_row_4, o_row_3, o_row_2, o_row_1, rtlc0n95: std_logic ;
   
   signal mem_wrn_current: std_logic_vector (2 DOWNTO 0) ;
   
   signal rtlc0n92, rtlcs0, not_rtlc0n196, rtlc0n196, not_rtlc0n207, 
      rtlc0n207, rtlc0n169, not_rtlcs0, not_first_bubble, rtlc0n225, 
      not_rtlc0n95, not_i_valid: std_logic ;
   
   signal mem_q_2_7_rename63: std_logic_vector (2 DOWNTO 1) ;
   
   signal mem_q_2_1_rename64: std_logic_vector (2 DOWNTO 2) ;
   
   signal mem_q_2_2_rename65: std_logic_vector (2 DOWNTO 2) ;
   
   signal mem_q_2_3_rename66: std_logic_vector (2 DOWNTO 2) ;
   
   signal mem_q_2_4_rename67: std_logic_vector (2 DOWNTO 2) ;
   
   signal mem_q_2_5_rename68: std_logic_vector (2 DOWNTO 2) ;
   
   signal mem_q_2_6_rename69: std_logic_vector (2 DOWNTO 2) ;
   
   signal mem_wrn: std_logic_vector (2 DOWNTO 0) ;
   
   signal mem_q_1_7_rename70: std_logic_vector (1 DOWNTO 0) ;
   
   signal mem_q_1_1_rename71: std_logic_vector (1 DOWNTO 1) ;
   
   signal mem_q_1_2_rename72: std_logic_vector (1 DOWNTO 1) ;
   
   signal mem_q_1_3_rename73: std_logic_vector (1 DOWNTO 1) ;
   
   signal mem_q_1_4_rename74: std_logic_vector (1 DOWNTO 1) ;
   
   signal mem_q_1_5_rename75: std_logic_vector (1 DOWNTO 1) ;
   
   signal mem_q_1_6_rename76: std_logic_vector (1 DOWNTO 1) ;
   
   signal mem_q_0_7_rename77: std_logic_vector (1 DOWNTO 0) ;
   
   signal mem_q_0_1_rename78: std_logic_vector (0 DOWNTO 0) ;
   
   signal mem_q_0_2_rename79: std_logic_vector (0 DOWNTO 0) ;
   
   signal mem_q_0_3_rename80: std_logic_vector (0 DOWNTO 0) ;
   
   signal mem_q_0_4_rename81: std_logic_vector (0 DOWNTO 0) ;
   
   signal mem_q_0_5_rename82: std_logic_vector (0 DOWNTO 0) ;
   
   signal mem_q_0_6_rename83: std_logic_vector (0 DOWNTO 0) ;
   
   signal mem_data: std_logic_vector (7 DOWNTO 0) ;
   
   signal o_column: std_logic_vector (7 DOWNTO 0) ;
   
   signal GND, PWR: std_logic ;
   
   signal DANGLING : std_logic_vector (15 downto 0 );

begin
   p_o_image1_9_7(1) <= o_image1_0_7_rename21(1) ;
   p_o_image1_9_1(0) <= o_image1_0_1_rename22(0) ;
   p_o_image1_9_2(0) <= o_image1_0_2_rename23(0) ;
   p_o_image1_9_3(0) <= o_image1_0_3_rename24(0) ;
   p_o_image1_9_4(0) <= o_image1_0_4_rename25(0) ;
   p_o_image1_9_5(0) <= o_image1_0_5_rename26(0) ;
   p_o_image1_9_6(0) <= o_image1_0_6_rename27(0) ;
   p_o_image1_9_7(0) <= o_image1_0_7_rename21(0) ;
   p_o_image1_8_7(1) <= o_image1_1_7_rename28(1) ;
   p_o_image1_8_1(1) <= o_image1_1_1_rename29(1) ;
   p_o_image1_8_2(1) <= o_image1_1_2_rename30(1) ;
   p_o_image1_8_3(1) <= o_image1_1_3_rename31(1) ;
   p_o_image1_8_4(1) <= o_image1_1_4_rename32(1) ;
   p_o_image1_8_5(1) <= o_image1_1_5_rename33(1) ;
   p_o_image1_8_6(1) <= o_image1_1_6_rename34(1) ;
   p_o_image1_8_7(0) <= o_image1_1_7_rename28(0) ;
   p_o_image1_7(2) <= o_image1_2_7_rename35(2) ;
   p_o_image1_1(2) <= o_image1_2_1_rename36(2) ;
   p_o_image1_2(2) <= o_image1_2_2_rename37(2) ;
   p_o_image1_3(2) <= o_image1_2_3_rename38(2) ;
   p_o_image1_4(2) <= o_image1_2_4_rename39(2) ;
   p_o_image1_5(2) <= o_image1_2_5_rename40(2) ;
   p_o_image1_6(2) <= o_image1_2_6_rename41(2) ;
   p_o_image1_7(1) <= o_image1_2_7_rename35(1) ;
   p_o_image2_9_7(1) <= o_image2_0_7_rename42(1) ;
   p_o_image2_9_1(0) <= o_image2_0_1_rename43(0) ;
   p_o_image2_9_2(0) <= o_image2_0_2_rename44(0) ;
   p_o_image2_9_3(0) <= o_image2_0_3_rename45(0) ;
   p_o_image2_9_4(0) <= o_image2_0_4_rename46(0) ;
   p_o_image2_9_5(0) <= o_image2_0_5_rename47(0) ;
   p_o_image2_9_6(0) <= o_image2_0_6_rename48(0) ;
   p_o_image2_9_7(0) <= o_image2_0_7_rename42(0) ;
   p_o_image2_8_7(1) <= o_image2_1_7_rename49(1) ;
   p_o_image2_8_1(1) <= o_image2_1_1_rename50(1) ;
   p_o_image2_8_2(1) <= o_image2_1_2_rename51(1) ;
   p_o_image2_8_3(1) <= o_image2_1_3_rename52(1) ;
   p_o_image2_8_4(1) <= o_image2_1_4_rename53(1) ;
   p_o_image2_8_5(1) <= o_image2_1_5_rename54(1) ;
   p_o_image2_8_6(1) <= o_image2_1_6_rename55(1) ;
   p_o_image2_8_7(0) <= o_image2_1_7_rename49(0) ;
   p_o_image2_7(2) <= o_image2_2_7_rename56(2) ;
   p_o_image2_1(2) <= o_image2_2_1_rename57(2) ;
   p_o_image2_2(2) <= o_image2_2_2_rename58(2) ;
   p_o_image2_3(2) <= o_image2_2_3_rename59(2) ;
   p_o_image2_4(2) <= o_image2_2_4_rename60(2) ;
   p_o_image2_5(2) <= o_image2_2_5_rename61(2) ;
   p_o_image2_6(2) <= o_image2_2_6_rename62(2) ;
   p_o_image2_7(1) <= o_image2_2_7_rename56(1) ;
   p_o_row(7) <= o_row_7 ;
   p_o_row(6) <= o_row_6 ;
   p_o_row(5) <= o_row_5 ;
   p_o_row(4) <= o_row_4 ;
   p_o_row(3) <= o_row_3 ;
   p_o_row(2) <= o_row_2 ;
   p_o_row(1) <= o_row_1 ;
   p_o_column(0) <= o_column(0) ;
   p_o_column(1) <= o_column(1) ;
   p_o_column(2) <= o_column(2) ;
   p_o_column(3) <= o_column(3) ;
   p_o_column(4) <= o_column(4) ;
   p_o_column(5) <= o_column(5) ;
   p_o_column(6) <= o_column(6) ;
   p_o_column(7) <= o_column(7) ;
   PWR <= '1' ;
   GND <= '0' ;
   u_mem1 : mem_8_8 port map ( address(7)=>o_column(7), address(6)=>
      o_column(6), address(5)=>o_column(5), address(4)=>o_column(4), 
      address(3)=>o_column(3), address(2)=>o_column(2), address(1)=>
      o_column(1), address(0)=>o_column(0), clock=>p_i_clock, data(7)=>
      mem_data(7), data(6)=>mem_data(6), data(5)=>mem_data(5), data(4)=>
      mem_data(4), data(3)=>mem_data(3), data(2)=>mem_data(2), data(1)=>
      mem_data(1), data(0)=>mem_data(0), wren=>mem_wrn(0), q(7)=>
      mem_q_0_7_rename77(0), q(6)=>mem_q_0_6_rename83(0), q(5)=>
      mem_q_0_5_rename82(0), q(4)=>mem_q_0_4_rename81(0), q(3)=>
      mem_q_0_3_rename80(0), q(2)=>mem_q_0_2_rename79(0), q(1)=>
      mem_q_0_1_rename78(0), q(0)=>mem_q_0_7_rename77(1));
   u_mem2 : mem_8_8 port map ( address(7)=>o_column(7), address(6)=>
      o_column(6), address(5)=>o_column(5), address(4)=>o_column(4), 
      address(3)=>o_column(3), address(2)=>o_column(2), address(1)=>
      o_column(1), address(0)=>o_column(0), clock=>p_i_clock, data(7)=>
      mem_data(7), data(6)=>mem_data(6), data(5)=>mem_data(5), data(4)=>
      mem_data(4), data(3)=>mem_data(3), data(2)=>mem_data(2), data(1)=>
      mem_data(1), data(0)=>mem_data(0), wren=>mem_wrn(1), q(7)=>
      mem_q_1_7_rename70(0), q(6)=>mem_q_1_6_rename76(1), q(5)=>
      mem_q_1_5_rename75(1), q(4)=>mem_q_1_4_rename74(1), q(3)=>
      mem_q_1_3_rename73(1), q(2)=>mem_q_1_2_rename72(1), q(1)=>
      mem_q_1_1_rename71(1), q(0)=>mem_q_1_7_rename70(1));
   u_mem3 : mem_8_8 port map ( address(7)=>o_column(7), address(6)=>
      o_column(6), address(5)=>o_column(5), address(4)=>o_column(4), 
      address(3)=>o_column(3), address(2)=>o_column(2), address(1)=>
      o_column(1), address(0)=>o_column(0), clock=>p_i_clock, data(7)=>
      mem_data(7), data(6)=>mem_data(6), data(5)=>mem_data(5), data(4)=>
      mem_data(4), data(3)=>mem_data(3), data(2)=>mem_data(2), data(1)=>
      mem_data(1), data(0)=>mem_data(0), wren=>mem_wrn(2), q(7)=>
      mem_q_2_7_rename63(1), q(6)=>mem_q_2_6_rename69(2), q(5)=>
      mem_q_2_5_rename68(2), q(4)=>mem_q_2_4_rename67(2), q(3)=>
      mem_q_2_3_rename66(2), q(2)=>mem_q_2_2_rename65(2), q(1)=>
      mem_q_2_1_rename64(2), q(0)=>mem_q_2_7_rename63(2));
   rtlc0n225 <= not_i_valid OR not_rtlc0n95 ;
   rtlc0n169 <= not_first_bubble OR not_rtlcs0 ;
   rtlc0n207 <= p_i_valid_rtlc_32_or_1(2) OR not_first_bubble ;
   not_rtlc0n207 <= NOT rtlc0n207 ;
   not_rtlc0n196 <= NOT rtlc0n196 ;
   not_rtlcs0 <= NOT rtlcs0 ;
   rtlc0n92 <= mem_wrn_current(0) OR mem_wrn_current(1) ;
   rtlc0n95 <= rtlc0n92 OR mem_wrn_current(2) ;
   not_rtlc0n95 <= NOT rtlc0n95 ;
   rtlc1_423_or_0 : or_7u_7u port map ( a(6)=>o_row_1, a(5)=>o_row_2, a(4)=>
      o_row_3, a(3)=>o_row_4, a(2)=>o_row_5, a(1)=>o_row_6, a(0)=>o_row_7, d
      =>rtlc1n272);
   rtlc_32_or_1 : or_3u_3u port map ( a(2)=>p_i_valid_rtlc_32_or_1(2), a(1)
      =>not_rtlcs0, a(0)=>not_first_bubble, d=>rtlc0n196);
   buffer2_select_1i1Bus7_0 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_7_rename77(1), b(1)
      =>buffer2_1n1ss1(0), b(0)=>mem_q_2_7_rename63(2), d=>buffer2_1n3ss1(0)
   );
   buffer2_select_1i1Bus7_1 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_1_rename78(0), b(1)
      =>buffer2_1n1ss1(1), b(0)=>mem_q_2_1_rename64(2), d=>buffer2_1n3ss1(1)
   );
   buffer2_select_1i1Bus7_2 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_2_rename79(0), b(1)
      =>buffer2_1n1ss1(2), b(0)=>mem_q_2_2_rename65(2), d=>buffer2_1n3ss1(2)
   );
   buffer2_select_1i1Bus7_3 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_3_rename80(0), b(1)
      =>buffer2_1n1ss1(3), b(0)=>mem_q_2_3_rename66(2), d=>buffer2_1n3ss1(3)
   );
   buffer2_select_1i1Bus7_4 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_4_rename81(0), b(1)
      =>buffer2_1n1ss1(4), b(0)=>mem_q_2_4_rename67(2), d=>buffer2_1n3ss1(4)
   );
   buffer2_select_1i1Bus7_5 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_5_rename82(0), b(1)
      =>buffer2_1n1ss1(5), b(0)=>mem_q_2_5_rename68(2), d=>buffer2_1n3ss1(5)
   );
   buffer2_select_1i1Bus7_6 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_6_rename83(0), b(1)
      =>buffer2_1n1ss1(6), b(0)=>mem_q_2_6_rename69(2), d=>buffer2_1n3ss1(6)
   );
   buffer2_select_1i1Bus7_7 : select_3_3 port map ( a(2)=>not_rtlcn225, a(1)
      =>mem_wrn_current(0), a(0)=>rtlcn97, b(2)=>mem_q_0_7_rename77(0), b(1)
      =>buffer2_1n1ss1(7), b(0)=>mem_q_2_7_rename63(1), d=>buffer2_1n3ss1(7)
   );
   buffer2_select_1i1Bus7_8 : select_3_3 port map ( a(2)=>not_rtlcn226, a(1)
      =>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_7_rename70(1), 
      b(1)=>buffer2_1n1ss1(0), b(0)=>mem_q_2_7_rename63(2), d=>
      buffer2_1n3ss1(8));
   buffer2_select_1i1Bus7_9 : select_3_3 port map ( a(2)=>not_rtlcn226, a(1)
      =>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_1_rename71(1), 
      b(1)=>buffer2_1n1ss1(1), b(0)=>mem_q_2_1_rename64(2), d=>
      buffer2_1n3ss1(9));
   buffer2_select_1i1Bus7_10 : select_3_3 port map ( a(2)=>not_rtlcn226, 
      a(1)=>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_2_rename72(1), 
      b(1)=>buffer2_1n1ss1(2), b(0)=>mem_q_2_2_rename65(2), d=>
      buffer2_1n3ss1(10));
   buffer2_select_1i1Bus7_11 : select_3_3 port map ( a(2)=>not_rtlcn226, 
      a(1)=>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_3_rename73(1), 
      b(1)=>buffer2_1n1ss1(3), b(0)=>mem_q_2_3_rename66(2), d=>
      buffer2_1n3ss1(11));
   buffer2_select_1i1Bus7_12 : select_3_3 port map ( a(2)=>not_rtlcn226, 
      a(1)=>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_4_rename74(1), 
      b(1)=>buffer2_1n1ss1(4), b(0)=>mem_q_2_4_rename67(2), d=>
      buffer2_1n3ss1(12));
   buffer2_select_1i1Bus7_13 : select_3_3 port map ( a(2)=>not_rtlcn226, 
      a(1)=>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_5_rename75(1), 
      b(1)=>buffer2_1n1ss1(5), b(0)=>mem_q_2_5_rename68(2), d=>
      buffer2_1n3ss1(13));
   buffer2_select_1i1Bus7_14 : select_3_3 port map ( a(2)=>not_rtlcn226, 
      a(1)=>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_6_rename76(1), 
      b(1)=>buffer2_1n1ss1(6), b(0)=>mem_q_2_6_rename69(2), d=>
      buffer2_1n3ss1(14));
   buffer2_select_1i1Bus7_15 : select_3_3 port map ( a(2)=>not_rtlcn226, 
      a(1)=>mem_wrn_current(1), a(0)=>rtlcn121, b(2)=>mem_q_1_7_rename70(0), 
      b(1)=>buffer2_1n1ss1(7), b(0)=>mem_q_2_7_rename63(1), d=>
      buffer2_1n3ss1(15));
   rtlcn97 <= rtlc1n272 AND mem_wrn_current(1) ;
   rtlcn121 <= rtlc1n272 AND mem_wrn_current(0) ;
   rtlcn217 <= mem_wrn_current(2) OR rtlc1n272 ;
   not_rtlcn225 <= NOT rtlcn225 ;
   not_rtlcn226 <= NOT rtlcn226 ;
   rtlc0n172 <= rtlc0n95 when p_i_valid_rtlc_32_or_1(2) = '1' else rtlc0n169
    ;
   buffer2_1n1ss1(0) <= mem_q_1_7_rename70(1) when rtlc1n272 = '1' else 
   mem_data(0) ;
   buffer2_1n1ss1(1) <= mem_q_1_1_rename71(1) when rtlc1n272 = '1' else 
   mem_data(1) ;
   buffer2_1n1ss1(2) <= mem_q_1_2_rename72(1) when rtlc1n272 = '1' else 
   mem_data(2) ;
   buffer2_1n1ss1(3) <= mem_q_1_3_rename73(1) when rtlc1n272 = '1' else 
   mem_data(3) ;
   buffer2_1n1ss1(4) <= mem_q_1_4_rename74(1) when rtlc1n272 = '1' else 
   mem_data(4) ;
   buffer2_1n1ss1(5) <= mem_q_1_5_rename75(1) when rtlc1n272 = '1' else 
   mem_data(5) ;
   buffer2_1n1ss1(6) <= mem_q_1_6_rename76(1) when rtlc1n272 = '1' else 
   mem_data(6) ;
   buffer2_1n1ss1(7) <= mem_q_1_7_rename70(0) when rtlc1n272 = '1' else 
   mem_data(7) ;
   buffer2_1n3ss1(16) <= mem_data(0) when rtlcn217 = '1' else 
   mem_q_2_7_rename63(2) ;
   buffer2_1n3ss1(17) <= mem_data(1) when rtlcn217 = '1' else 
   mem_q_2_1_rename64(2) ;
   buffer2_1n3ss1(18) <= mem_data(2) when rtlcn217 = '1' else 
   mem_q_2_2_rename65(2) ;
   buffer2_1n3ss1(19) <= mem_data(3) when rtlcn217 = '1' else 
   mem_q_2_3_rename66(2) ;
   buffer2_1n3ss1(20) <= mem_data(4) when rtlcn217 = '1' else 
   mem_q_2_4_rename67(2) ;
   buffer2_1n3ss1(21) <= mem_data(5) when rtlcn217 = '1' else 
   mem_q_2_5_rename68(2) ;
   buffer2_1n3ss1(22) <= mem_data(6) when rtlcn217 = '1' else 
   mem_q_2_6_rename69(2) ;
   buffer2_1n3ss1(23) <= mem_data(7) when rtlcn217 = '1' else 
   mem_q_2_7_rename63(1) ;
   not_rtlc0n172 <= NOT rtlc0n172 ;
   not_first_bubble <= NOT first_bubble ;
   not_i_valid <= NOT p_i_valid_rtlc_32_or_1(2) ;
   rtlc_522_and_18 : and_8u_8u port map ( a(7)=>o_column(7), a(6)=>
      o_column(6), a(5)=>o_column(5), a(4)=>o_column(4), a(3)=>o_column(3), 
      a(2)=>o_column(2), a(1)=>o_column(1), a(0)=>o_column(0), d=>rtlcs0);
   mem_wrn_current_0n4ss1(1) <= mem_wrn_current(0) AND not_i_valid ;
   mem_wrn_current_0n4ss1(2) <= mem_wrn_current(1) AND not_i_valid ;
   mem_wrn_current_0n4ss1(0) <= mem_wrn_current(2) OR 
   p_i_valid_rtlc_32_or_1(2) ;
   rtlcn225 <= mem_wrn_current(0) OR rtlcn97 ;
   rtlcn226 <= mem_wrn_current(1) OR rtlcn121 ;
   modgen_counter_o_row : counter_up_cnt_en_clock_0_8 port map ( clock=>
      p_i_clock, q(7)=>o_row_7, q(6)=>o_row_6, q(5)=>o_row_5, q(4)=>o_row_4, 
      q(3)=>o_row_3, q(2)=>o_row_2, q(1)=>o_row_1, q(0)=>p_o_row(0), clk_en
      =>PWR, aclear=>GND, sload=>GND, data(7)=>DANGLING(0), data(6)=>
      DANGLING(1), data(5)=>DANGLING(2), data(4)=>DANGLING(3), data(3)=>
      DANGLING(4), data(2)=>DANGLING(5), data(1)=>DANGLING(6), data(0)=>
      DANGLING(7), aset=>GND, sclear=>GND, updn=>PWR, cnt_en=>not_rtlc0n196
   );
   modgen_counter_o_column : counter_up_sclear_clock_clk_en_0_8 port map ( 
      clock=>p_i_clock, q(7)=>o_column(7), q(6)=>o_column(6), q(5)=>
      o_column(5), q(4)=>o_column(4), q(3)=>o_column(3), q(2)=>o_column(2), 
      q(1)=>o_column(1), q(0)=>o_column(0), clk_en=>not_rtlc0n207, aclear=>
      GND, sload=>GND, data(7)=>DANGLING(8), data(6)=>DANGLING(9), data(5)=>
      DANGLING(10), data(4)=>DANGLING(11), data(3)=>DANGLING(12), data(2)=>
      DANGLING(13), data(1)=>DANGLING(14), data(0)=>DANGLING(15), aset=>GND, 
      sclear=>rtlcs0, updn=>PWR, cnt_en=>PWR);
   not_rtlc0n225 <= NOT rtlc0n225 ;
   rtlcn229 <= mem_wrn_current(2) AND not_rtlc0n225 ;
   rtlcn231 <= mem_wrn_current(1) AND not_rtlc0n225 ;
   rtlcn233 <= mem_wrn_current(0) OR not_rtlc0n95 ;
   rtlcn234 <= rtlcn233 AND p_i_valid_rtlc_32_or_1(2) ;
   DFFPCE (mem_wrn_current_0n4ss1(2),GND,GND,not_rtlc0n172,p_i_clock,
   mem_wrn_current(2)) ;
   DFFPCE (mem_wrn_current_0n4ss1(1),GND,GND,not_rtlc0n172,p_i_clock,
   mem_wrn_current(1)) ;
   DFFPCE (mem_wrn_current_0n4ss1(0),GND,GND,not_rtlc0n172,p_i_clock,
   mem_wrn_current(0)) ;
   DFFPCE (p_i_pixel(7),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(7)) ;
   DFFPCE (p_i_pixel(6),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(6)) ;
   DFFPCE (p_i_pixel(5),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(5)) ;
   DFFPCE (p_i_pixel(4),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(4)) ;
   DFFPCE (p_i_pixel(3),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(3)) ;
   DFFPCE (p_i_pixel(2),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(2)) ;
   DFFPCE (p_i_pixel(1),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(1)) ;
   DFFPCE (p_i_pixel(0),GND,GND,p_i_valid_rtlc_32_or_1(2),p_i_clock,
   mem_data(0)) ;
   DFFPCE (buffer2_1n3ss1(23),GND,GND,first_bubble,p_i_clock,
   o_image2_2_7_rename56(1)) ;
   DFFPCE (buffer2_1n3ss1(22),GND,GND,first_bubble,p_i_clock,
   o_image2_2_6_rename62(2)) ;
   DFFPCE (buffer2_1n3ss1(21),GND,GND,first_bubble,p_i_clock,
   o_image2_2_5_rename61(2)) ;
   DFFPCE (buffer2_1n3ss1(20),GND,GND,first_bubble,p_i_clock,
   o_image2_2_4_rename60(2)) ;
   DFFPCE (buffer2_1n3ss1(19),GND,GND,first_bubble,p_i_clock,
   o_image2_2_3_rename59(2)) ;
   DFFPCE (buffer2_1n3ss1(18),GND,GND,first_bubble,p_i_clock,
   o_image2_2_2_rename58(2)) ;
   DFFPCE (buffer2_1n3ss1(17),GND,GND,first_bubble,p_i_clock,
   o_image2_2_1_rename57(2)) ;
   DFFPCE (buffer2_1n3ss1(16),GND,GND,first_bubble,p_i_clock,
   o_image2_2_7_rename56(2)) ;
   DFFPCE (buffer2_1n3ss1(15),GND,GND,first_bubble,p_i_clock,
   o_image2_1_7_rename49(0)) ;
   DFFPCE (buffer2_1n3ss1(14),GND,GND,first_bubble,p_i_clock,
   o_image2_1_6_rename55(1)) ;
   DFFPCE (buffer2_1n3ss1(13),GND,GND,first_bubble,p_i_clock,
   o_image2_1_5_rename54(1)) ;
   DFFPCE (buffer2_1n3ss1(12),GND,GND,first_bubble,p_i_clock,
   o_image2_1_4_rename53(1)) ;
   DFFPCE (buffer2_1n3ss1(11),GND,GND,first_bubble,p_i_clock,
   o_image2_1_3_rename52(1)) ;
   DFFPCE (buffer2_1n3ss1(10),GND,GND,first_bubble,p_i_clock,
   o_image2_1_2_rename51(1)) ;
   DFFPCE (buffer2_1n3ss1(9),GND,GND,first_bubble,p_i_clock,
   o_image2_1_1_rename50(1)) ;
   DFFPCE (buffer2_1n3ss1(8),GND,GND,first_bubble,p_i_clock,
   o_image2_1_7_rename49(1)) ;
   DFFPCE (buffer2_1n3ss1(7),GND,GND,first_bubble,p_i_clock,
   o_image2_0_7_rename42(0)) ;
   DFFPCE (buffer2_1n3ss1(6),GND,GND,first_bubble,p_i_clock,
   o_image2_0_6_rename48(0)) ;
   DFFPCE (buffer2_1n3ss1(5),GND,GND,first_bubble,p_i_clock,
   o_image2_0_5_rename47(0)) ;
   DFFPCE (buffer2_1n3ss1(4),GND,GND,first_bubble,p_i_clock,
   o_image2_0_4_rename46(0)) ;
   DFFPCE (buffer2_1n3ss1(3),GND,GND,first_bubble,p_i_clock,
   o_image2_0_3_rename45(0)) ;
   DFFPCE (buffer2_1n3ss1(2),GND,GND,first_bubble,p_i_clock,
   o_image2_0_2_rename44(0)) ;
   DFFPCE (buffer2_1n3ss1(1),GND,GND,first_bubble,p_i_clock,
   o_image2_0_1_rename43(0)) ;
   DFFPCE (buffer2_1n3ss1(0),GND,GND,first_bubble,p_i_clock,
   o_image2_0_7_rename42(1)) ;
   DFFPCE (o_image2_2_7_rename56(1),GND,GND,first_bubble,p_i_clock,
   o_image1_2_7_rename35(1)) ;
   DFFPCE (o_image2_2_6_rename62(2),GND,GND,first_bubble,p_i_clock,
   o_image1_2_6_rename41(2)) ;
   DFFPCE (o_image2_2_5_rename61(2),GND,GND,first_bubble,p_i_clock,
   o_image1_2_5_rename40(2)) ;
   DFFPCE (o_image2_2_4_rename60(2),GND,GND,first_bubble,p_i_clock,
   o_image1_2_4_rename39(2)) ;
   DFFPCE (o_image2_2_3_rename59(2),GND,GND,first_bubble,p_i_clock,
   o_image1_2_3_rename38(2)) ;
   DFFPCE (o_image2_2_2_rename58(2),GND,GND,first_bubble,p_i_clock,
   o_image1_2_2_rename37(2)) ;
   DFFPCE (o_image2_2_1_rename57(2),GND,GND,first_bubble,p_i_clock,
   o_image1_2_1_rename36(2)) ;
   DFFPCE (o_image2_2_7_rename56(2),GND,GND,first_bubble,p_i_clock,
   o_image1_2_7_rename35(2)) ;
   DFFPCE (o_image2_1_7_rename49(0),GND,GND,first_bubble,p_i_clock,
   o_image1_1_7_rename28(0)) ;
   DFFPCE (o_image2_1_6_rename55(1),GND,GND,first_bubble,p_i_clock,
   o_image1_1_6_rename34(1)) ;
   DFFPCE (o_image2_1_5_rename54(1),GND,GND,first_bubble,p_i_clock,
   o_image1_1_5_rename33(1)) ;
   DFFPCE (o_image2_1_4_rename53(1),GND,GND,first_bubble,p_i_clock,
   o_image1_1_4_rename32(1)) ;
   DFFPCE (o_image2_1_3_rename52(1),GND,GND,first_bubble,p_i_clock,
   o_image1_1_3_rename31(1)) ;
   DFFPCE (o_image2_1_2_rename51(1),GND,GND,first_bubble,p_i_clock,
   o_image1_1_2_rename30(1)) ;
   DFFPCE (o_image2_1_1_rename50(1),GND,GND,first_bubble,p_i_clock,
   o_image1_1_1_rename29(1)) ;
   DFFPCE (o_image2_1_7_rename49(1),GND,GND,first_bubble,p_i_clock,
   o_image1_1_7_rename28(1)) ;
   DFFPCE (o_image2_0_7_rename42(0),GND,GND,first_bubble,p_i_clock,
   o_image1_0_7_rename21(0)) ;
   DFFPCE (o_image2_0_6_rename48(0),GND,GND,first_bubble,p_i_clock,
   o_image1_0_6_rename27(0)) ;
   DFFPCE (o_image2_0_5_rename47(0),GND,GND,first_bubble,p_i_clock,
   o_image1_0_5_rename26(0)) ;
   DFFPCE (o_image2_0_4_rename46(0),GND,GND,first_bubble,p_i_clock,
   o_image1_0_4_rename25(0)) ;
   DFFPCE (o_image2_0_3_rename45(0),GND,GND,first_bubble,p_i_clock,
   o_image1_0_3_rename24(0)) ;
   DFFPCE (o_image2_0_2_rename44(0),GND,GND,first_bubble,p_i_clock,
   o_image1_0_2_rename23(0)) ;
   DFFPCE (o_image2_0_1_rename43(0),GND,GND,first_bubble,p_i_clock,
   o_image1_0_1_rename22(0)) ;
   DFFPCE (o_image2_0_7_rename42(1),GND,GND,first_bubble,p_i_clock,
   o_image1_0_7_rename21(1)) ;
   DFFPCE (o_image1_2_7_rename35(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_7(1)) ;
   DFFPCE (o_image1_2_6_rename41(2),GND,GND,first_bubble,p_i_clock,
   p_o_image0_6(2)) ;
   DFFPCE (o_image1_2_5_rename40(2),GND,GND,first_bubble,p_i_clock,
   p_o_image0_5(2)) ;
   DFFPCE (o_image1_2_4_rename39(2),GND,GND,first_bubble,p_i_clock,
   p_o_image0_4(2)) ;
   DFFPCE (o_image1_2_3_rename38(2),GND,GND,first_bubble,p_i_clock,
   p_o_image0_3(2)) ;
   DFFPCE (o_image1_2_2_rename37(2),GND,GND,first_bubble,p_i_clock,
   p_o_image0_2(2)) ;
   DFFPCE (o_image1_2_1_rename36(2),GND,GND,first_bubble,p_i_clock,
   p_o_image0_1(2)) ;
   DFFPCE (o_image1_2_7_rename35(2),GND,GND,first_bubble,p_i_clock,
   p_o_image0_7(2)) ;
   DFFPCE (o_image1_1_7_rename28(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_7(0)) ;
   DFFPCE (o_image1_1_6_rename34(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_6(1)) ;
   DFFPCE (o_image1_1_5_rename33(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_5(1)) ;
   DFFPCE (o_image1_1_4_rename32(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_4(1)) ;
   DFFPCE (o_image1_1_3_rename31(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_3(1)) ;
   DFFPCE (o_image1_1_2_rename30(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_2(1)) ;
   DFFPCE (o_image1_1_1_rename29(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_1(1)) ;
   DFFPCE (o_image1_1_7_rename28(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_8_7(1)) ;
   DFFPCE (o_image1_0_7_rename21(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_7(0)) ;
   DFFPCE (o_image1_0_6_rename27(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_6(0)) ;
   DFFPCE (o_image1_0_5_rename26(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_5(0)) ;
   DFFPCE (o_image1_0_4_rename25(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_4(0)) ;
   DFFPCE (o_image1_0_3_rename24(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_3(0)) ;
   DFFPCE (o_image1_0_2_rename23(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_2(0)) ;
   DFFPCE (o_image1_0_1_rename22(0),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_1(0)) ;
   DFFPCE (o_image1_0_7_rename21(1),GND,GND,first_bubble,p_i_clock,
   p_o_image0_9_7(1)) ;
   DFFPC (rtlcn229,GND,GND,p_i_clock,mem_wrn(2)) ;
   DFFPC (rtlcn231,GND,GND,p_i_clock,mem_wrn(1)) ;
   DFFPC (rtlcn234,GND,GND,p_i_clock,mem_wrn(0)) ;
   DFFPC (p_i_valid_rtlc_32_or_1(2),GND,GND,p_i_clock,first_bubble) ;
end main_unfold_1492 ;

library IEEE;library altera_mf;library lpm;library altera; 
 use IEEE.STD_LOGIC_1164.ALL;
 use altera_mf.altera_mf_components.all, lpm.lpm_components.all, altera.altera_primitives_components.all;

entity kirsch is 
   port (
      i_clock : IN std_logic ;
      i_reset : IN std_logic ;
      i_valid : IN std_logic ;
      i_pixel : IN std_logic_vector (7 DOWNTO 0) ;
      o_valid : OUT std_logic ;
      o_edge : OUT std_logic ;
      o_dir : OUT std_logic_vector (2 DOWNTO 0) ;
      o_mode : OUT std_logic_vector (1 DOWNTO 0) ;
      o_row : OUT std_logic_vector (7 DOWNTO 0) ;
      o_pixel : OUT std_logic_vector (7 DOWNTO 0) ;
      o_column : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image0_0 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image0_1 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image0_2 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image1_0 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image1_1 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image1_2 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image2_0 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image2_1 : OUT std_logic_vector (7 DOWNTO 0) ;
      o_image2_2 : OUT std_logic_vector (7 DOWNTO 0) ;
      debug_key : IN std_logic_vector (3 DOWNTO 1) ;
      debug_switch : IN std_logic_vector (17 DOWNTO 0) ;
      debug_led_red : OUT std_logic_vector (17 DOWNTO 0) ;
      debug_led_grn : OUT std_logic_vector (5 DOWNTO 0) ;
      debug_num_0 : OUT std_logic_vector (3 DOWNTO 0) ;
      debug_num_1 : OUT std_logic_vector (3 DOWNTO 0) ;
      debug_num_2 : OUT std_logic_vector (3 DOWNTO 0) ;
      debug_num_3 : OUT std_logic_vector (3 DOWNTO 0) ;
      debug_num_4 : OUT std_logic_vector (3 DOWNTO 0) ;
      debug_num_5 : OUT std_logic_vector (3 DOWNTO 0)) ;
end kirsch ;

architecture main of kirsch is 
   component memory_notri
      port (
         p_o_image0_9_7 : OUT std_logic_vector (1 DOWNTO 0) ;
         p_o_image0_9_1 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image0_9_2 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image0_9_3 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image0_9_4 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image0_9_5 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image0_9_6 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image0_8_7 : OUT std_logic_vector (1 DOWNTO 0) ;
         p_o_image0_8_1 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image0_8_2 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image0_8_3 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image0_8_4 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image0_8_5 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image0_8_6 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image0_7 : OUT std_logic_vector (2 DOWNTO 1) ;
         p_o_image0_1 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image0_2 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image0_3 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image0_4 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image0_5 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image0_6 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image1_9_7 : OUT std_logic_vector (1 DOWNTO 0) ;
         p_o_image1_9_1 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image1_9_2 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image1_9_3 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image1_9_4 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image1_9_5 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image1_9_6 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image1_8_7 : OUT std_logic_vector (1 DOWNTO 0) ;
         p_o_image1_8_1 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image1_8_2 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image1_8_3 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image1_8_4 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image1_8_5 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image1_8_6 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image1_7 : OUT std_logic_vector (2 DOWNTO 1) ;
         p_o_image1_1 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image1_2 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image1_3 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image1_4 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image1_5 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image1_6 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image2_9_7 : OUT std_logic_vector (1 DOWNTO 0) ;
         p_o_image2_9_1 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image2_9_2 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image2_9_3 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image2_9_4 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image2_9_5 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image2_9_6 : OUT std_logic_vector (0 DOWNTO 0) ;
         p_o_image2_8_7 : OUT std_logic_vector (1 DOWNTO 0) ;
         p_o_image2_8_1 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image2_8_2 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image2_8_3 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image2_8_4 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image2_8_5 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image2_8_6 : OUT std_logic_vector (1 DOWNTO 1) ;
         p_o_image2_7 : OUT std_logic_vector (2 DOWNTO 1) ;
         p_o_image2_1 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image2_2 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image2_3 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image2_4 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image2_5 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_o_image2_6 : OUT std_logic_vector (2 DOWNTO 2) ;
         p_i_pixel : IN std_logic_vector (7 DOWNTO 0) ;
         p_o_row : OUT std_logic_vector (7 DOWNTO 0) ;
         p_i_valid_rtlc_32_or_1 : IN std_logic_vector (2 DOWNTO 2) ;
         p_i_clock : IN std_logic ;
         p_o_column : OUT std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   signal debug_num_5_1_EXMPLR249, debug_num_5_0_EXMPLR250: std_logic ;

begin
   debug_led_red(17) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(16) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(15) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(14) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(13) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(12) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(11) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(10) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(9) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(8) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(7) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(6) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(5) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(4) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(3) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(2) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(1) <= debug_num_5_0_EXMPLR250 ;
   debug_led_red(0) <= debug_num_5_0_EXMPLR250 ;
   debug_led_grn(5) <= debug_num_5_0_EXMPLR250 ;
   debug_led_grn(4) <= debug_num_5_0_EXMPLR250 ;
   debug_led_grn(3) <= debug_num_5_0_EXMPLR250 ;
   debug_led_grn(2) <= debug_num_5_0_EXMPLR250 ;
   debug_led_grn(1) <= debug_num_5_0_EXMPLR250 ;
   debug_led_grn(0) <= debug_num_5_0_EXMPLR250 ;
   debug_num_0(3) <= debug_num_5_0_EXMPLR250 ;
   debug_num_0(2) <= debug_num_5_1_EXMPLR249 ;
   debug_num_0(1) <= debug_num_5_1_EXMPLR249 ;
   debug_num_0(0) <= debug_num_5_1_EXMPLR249 ;
   debug_num_1(3) <= debug_num_5_0_EXMPLR250 ;
   debug_num_1(2) <= debug_num_5_0_EXMPLR250 ;
   debug_num_1(1) <= debug_num_5_1_EXMPLR249 ;
   debug_num_1(0) <= debug_num_5_0_EXMPLR250 ;
   debug_num_2(3) <= debug_num_5_0_EXMPLR250 ;
   debug_num_2(2) <= debug_num_5_0_EXMPLR250 ;
   debug_num_2(1) <= debug_num_5_1_EXMPLR249 ;
   debug_num_2(0) <= debug_num_5_1_EXMPLR249 ;
   debug_num_3(3) <= debug_num_5_1_EXMPLR249 ;
   debug_num_3(2) <= debug_num_5_1_EXMPLR249 ;
   debug_num_3(1) <= debug_num_5_1_EXMPLR249 ;
   debug_num_3(0) <= debug_num_5_0_EXMPLR250 ;
   debug_num_4(3) <= debug_num_5_1_EXMPLR249 ;
   debug_num_4(2) <= debug_num_5_1_EXMPLR249 ;
   debug_num_4(1) <= debug_num_5_0_EXMPLR250 ;
   debug_num_4(0) <= debug_num_5_0_EXMPLR250 ;
   debug_num_5(3) <= debug_num_5_1_EXMPLR249 ;
   debug_num_5(2) <= debug_num_5_1_EXMPLR249 ;
   debug_num_5(1) <= debug_num_5_1_EXMPLR249 ;
   debug_num_5(0) <= debug_num_5_0_EXMPLR250 ;
   debug_num_5_1_EXMPLR249 <= '1' ;
   debug_num_5_0_EXMPLR250 <= '0' ;
   o_valid <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_edge <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_dir(0) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_dir(1) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_dir(2) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_mode(0) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_mode(1) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(0) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(1) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(2) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(3) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(4) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(5) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(6) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   o_pixel(7) <= debug_num_5_0_EXMPLR250 when debug_num_5_0_EXMPLR250
    = '1' else 'Z' ;
   u_memory : memory_notri port map ( p_o_image0_9_7(1)=>o_image0_0(0), 
      p_o_image0_9_7(0)=>o_image0_0(7), p_o_image0_9_1(0)=>o_image0_0(1), 
      p_o_image0_9_2(0)=>o_image0_0(2), p_o_image0_9_3(0)=>o_image0_0(3), 
      p_o_image0_9_4(0)=>o_image0_0(4), p_o_image0_9_5(0)=>o_image0_0(5), 
      p_o_image0_9_6(0)=>o_image0_0(6), p_o_image0_8_7(1)=>o_image0_1(0), 
      p_o_image0_8_7(0)=>o_image0_1(7), p_o_image0_8_1(1)=>o_image0_1(1), 
      p_o_image0_8_2(1)=>o_image0_1(2), p_o_image0_8_3(1)=>o_image0_1(3), 
      p_o_image0_8_4(1)=>o_image0_1(4), p_o_image0_8_5(1)=>o_image0_1(5), 
      p_o_image0_8_6(1)=>o_image0_1(6), p_o_image0_7(2)=>o_image0_2(0), 
      p_o_image0_7(1)=>o_image0_2(7), p_o_image0_1(2)=>o_image0_2(1), 
      p_o_image0_2(2)=>o_image0_2(2), p_o_image0_3(2)=>o_image0_2(3), 
      p_o_image0_4(2)=>o_image0_2(4), p_o_image0_5(2)=>o_image0_2(5), 
      p_o_image0_6(2)=>o_image0_2(6), p_o_image1_9_7(1)=>o_image1_0(0), 
      p_o_image1_9_7(0)=>o_image1_0(7), p_o_image1_9_1(0)=>o_image1_0(1), 
      p_o_image1_9_2(0)=>o_image1_0(2), p_o_image1_9_3(0)=>o_image1_0(3), 
      p_o_image1_9_4(0)=>o_image1_0(4), p_o_image1_9_5(0)=>o_image1_0(5), 
      p_o_image1_9_6(0)=>o_image1_0(6), p_o_image1_8_7(1)=>o_image1_1(0), 
      p_o_image1_8_7(0)=>o_image1_1(7), p_o_image1_8_1(1)=>o_image1_1(1), 
      p_o_image1_8_2(1)=>o_image1_1(2), p_o_image1_8_3(1)=>o_image1_1(3), 
      p_o_image1_8_4(1)=>o_image1_1(4), p_o_image1_8_5(1)=>o_image1_1(5), 
      p_o_image1_8_6(1)=>o_image1_1(6), p_o_image1_7(2)=>o_image1_2(0), 
      p_o_image1_7(1)=>o_image1_2(7), p_o_image1_1(2)=>o_image1_2(1), 
      p_o_image1_2(2)=>o_image1_2(2), p_o_image1_3(2)=>o_image1_2(3), 
      p_o_image1_4(2)=>o_image1_2(4), p_o_image1_5(2)=>o_image1_2(5), 
      p_o_image1_6(2)=>o_image1_2(6), p_o_image2_9_7(1)=>o_image2_0(0), 
      p_o_image2_9_7(0)=>o_image2_0(7), p_o_image2_9_1(0)=>o_image2_0(1), 
      p_o_image2_9_2(0)=>o_image2_0(2), p_o_image2_9_3(0)=>o_image2_0(3), 
      p_o_image2_9_4(0)=>o_image2_0(4), p_o_image2_9_5(0)=>o_image2_0(5), 
      p_o_image2_9_6(0)=>o_image2_0(6), p_o_image2_8_7(1)=>o_image2_1(0), 
      p_o_image2_8_7(0)=>o_image2_1(7), p_o_image2_8_1(1)=>o_image2_1(1), 
      p_o_image2_8_2(1)=>o_image2_1(2), p_o_image2_8_3(1)=>o_image2_1(3), 
      p_o_image2_8_4(1)=>o_image2_1(4), p_o_image2_8_5(1)=>o_image2_1(5), 
      p_o_image2_8_6(1)=>o_image2_1(6), p_o_image2_7(2)=>o_image2_2(0), 
      p_o_image2_7(1)=>o_image2_2(7), p_o_image2_1(2)=>o_image2_2(1), 
      p_o_image2_2(2)=>o_image2_2(2), p_o_image2_3(2)=>o_image2_2(3), 
      p_o_image2_4(2)=>o_image2_2(4), p_o_image2_5(2)=>o_image2_2(5), 
      p_o_image2_6(2)=>o_image2_2(6), p_i_pixel(7)=>i_pixel(7), p_i_pixel(6)
      =>i_pixel(6), p_i_pixel(5)=>i_pixel(5), p_i_pixel(4)=>i_pixel(4), 
      p_i_pixel(3)=>i_pixel(3), p_i_pixel(2)=>i_pixel(2), p_i_pixel(1)=>
      i_pixel(1), p_i_pixel(0)=>i_pixel(0), p_o_row(7)=>o_row(7), p_o_row(6)
      =>o_row(6), p_o_row(5)=>o_row(5), p_o_row(4)=>o_row(4), p_o_row(3)=>
      o_row(3), p_o_row(2)=>o_row(2), p_o_row(1)=>o_row(1), p_o_row(0)=>
      o_row(0), p_i_valid_rtlc_32_or_1(2)=>i_valid, p_i_clock=>i_clock, 
      p_o_column(7)=>o_column(7), p_o_column(6)=>o_column(6), p_o_column(5)
      =>o_column(5), p_o_column(4)=>o_column(4), p_o_column(3)=>o_column(3), 
      p_o_column(2)=>o_column(2), p_o_column(1)=>o_column(1), p_o_column(0)
      =>o_column(0));
end main ;

