library verilog;
use verilog.vl_types.all;
entity flow_notri is
    port(
        p_i_valid_ix261 : in     vl_logic_vector(0 downto 0);
        p_i_mode        : in     vl_logic_vector(1 downto 0);
        p_o_row         : out    vl_logic_vector(7 downto 0);
        p_i_row         : in     vl_logic_vector(7 downto 0);
        p_o_valid       : out    vl_logic;
        p_debug_valid   : out    vl_logic;
        p_i_clock       : in     vl_logic;
        p_i2            : in     vl_logic_vector(7 downto 0);
        p_i1            : in     vl_logic_vector(7 downto 0);
        p_b3            : in     vl_logic_vector(7 downto 0);
        p_b2            : in     vl_logic_vector(7 downto 0);
        p_b1            : in     vl_logic_vector(7 downto 0);
        p_t3            : in     vl_logic_vector(7 downto 0);
        p_t2            : in     vl_logic_vector(7 downto 0);
        p_t1            : in     vl_logic_vector(7 downto 0);
        p_o_mode        : out    vl_logic_vector(1 downto 0);
        p_o_dir         : out    vl_logic_vector(2 downto 0);
        p_o_edge        : out    vl_logic;
        p_debug_num_6   : out    vl_logic;
        p_debug_num_7   : out    vl_logic;
        p_debug_num_3   : out    vl_logic_vector(12 downto 0);
        p_debug_num_4   : out    vl_logic_vector(12 downto 0);
        p_i_reset       : in     vl_logic;
        p_debug_num_2   : out    vl_logic_vector(12 downto 0);
        p_debug_num_1   : out    vl_logic_vector(10 downto 0);
        p_debug_num_0   : out    vl_logic_vector(12 downto 0);
        p_ix259_ix248_nx13: out    vl_logic;
        p_ix259_ix249_nx13: out    vl_logic;
        p_ix259_ix250_nx13: out    vl_logic;
        p_ix259_ix251_nx13: out    vl_logic;
        p_ix259_ix252_nx13: out    vl_logic;
        p_ix259_ix253_nx13: out    vl_logic;
        p_ix259_ix254_nx13: out    vl_logic;
        p_ix259_ix255_nx13: out    vl_logic;
        p_not_rtlc5n47  : out    vl_logic;
        \p_p23_10_\     : out    vl_logic;
        \p_p23_9_\      : out    vl_logic;
        \p_p23_8_\      : out    vl_logic;
        \p_p23_7_\      : out    vl_logic;
        \p_p23_6_\      : out    vl_logic;
        \p_p23_5_\      : out    vl_logic;
        \p_p23_4_\      : out    vl_logic;
        \p_p23_3_\      : out    vl_logic;
        \p_p23_2_\      : out    vl_logic;
        \p_p23_1_\      : out    vl_logic;
        \p_p23_0_\      : out    vl_logic;
        \p_p21_4n0r2_12_\: out    vl_logic;
        \p_p21_4n0r2_11_\: out    vl_logic;
        \p_p21_4n0r2_10_\: out    vl_logic;
        \p_p21_4n0r2_9_\: out    vl_logic;
        \p_p21_4n0r2_8_\: out    vl_logic;
        \p_p21_4n0r2_7_\: out    vl_logic;
        \p_p21_4n0r2_6_\: out    vl_logic;
        \p_p21_4n0r2_5_\: out    vl_logic;
        \p_p21_4n0r2_4_\: out    vl_logic;
        \p_p21_4n0r2_3_\: out    vl_logic;
        \p_p21_4n0r2_2_\: out    vl_logic;
        \p_p21_4n0r2_1_\: out    vl_logic;
        \p_p21_4n0r3_0_\: out    vl_logic;
        \p_p22_4n0r2_12_\: out    vl_logic;
        \p_p22_4n0r2_11_\: out    vl_logic;
        \p_p22_4n0r2_10_\: out    vl_logic;
        \p_p22_4n0r2_9_\: out    vl_logic;
        \p_p22_4n0r2_8_\: out    vl_logic;
        \p_p22_4n0r2_7_\: out    vl_logic;
        \p_p22_4n0r2_6_\: out    vl_logic;
        \p_p22_4n0r2_5_\: out    vl_logic;
        \p_p22_4n0r2_4_\: out    vl_logic;
        \p_p22_4n0r2_3_\: out    vl_logic;
        \p_p22_4n0r2_2_\: out    vl_logic;
        \p_p22_4n0r2_1_\: out    vl_logic;
        \p_p22_4n0r3_0_\: out    vl_logic;
        \p_p5m_1_\      : out    vl_logic;
        \p_p5m_0_\      : out    vl_logic
    );
end flow_notri;
