library verilog;
use verilog.vl_types.all;
entity memory_notri is
    port(
        p_i_pixel       : in     vl_logic_vector(7 downto 0);
        p_o_row         : out    vl_logic_vector(7 downto 0);
        p_o_valid       : out    vl_logic;
        p_o_image0_9_7  : out    vl_logic_vector(1 downto 0);
        p_o_image0_9_1  : out    vl_logic_vector(0 downto 0);
        p_o_image0_9_2  : out    vl_logic_vector(0 downto 0);
        p_o_image0_9_3  : out    vl_logic_vector(0 downto 0);
        p_o_image0_9_4  : out    vl_logic_vector(0 downto 0);
        p_o_image0_9_5  : out    vl_logic_vector(0 downto 0);
        p_o_image0_9_6  : out    vl_logic_vector(0 downto 0);
        p_o_image0_8_7  : out    vl_logic_vector(1 downto 0);
        p_o_image0_8_1  : out    vl_logic_vector(1 downto 1);
        p_o_image0_8_2  : out    vl_logic_vector(1 downto 1);
        p_o_image0_8_3  : out    vl_logic_vector(1 downto 1);
        p_o_image0_8_4  : out    vl_logic_vector(1 downto 1);
        p_o_image0_8_5  : out    vl_logic_vector(1 downto 1);
        p_o_image0_8_6  : out    vl_logic_vector(1 downto 1);
        p_o_image0_7    : out    vl_logic_vector(2 downto 1);
        p_o_image0_1    : out    vl_logic_vector(2 downto 2);
        p_o_image0_2    : out    vl_logic_vector(2 downto 2);
        p_o_image0_3    : out    vl_logic_vector(2 downto 2);
        p_o_image0_4    : out    vl_logic_vector(2 downto 2);
        p_o_image0_5    : out    vl_logic_vector(2 downto 2);
        p_o_image0_6    : out    vl_logic_vector(2 downto 2);
        p_o_image1_9_7  : out    vl_logic_vector(1 downto 0);
        p_o_image1_9_1  : out    vl_logic_vector(0 downto 0);
        p_o_image1_9_2  : out    vl_logic_vector(0 downto 0);
        p_o_image1_9_3  : out    vl_logic_vector(0 downto 0);
        p_o_image1_9_4  : out    vl_logic_vector(0 downto 0);
        p_o_image1_9_5  : out    vl_logic_vector(0 downto 0);
        p_o_image1_9_6  : out    vl_logic_vector(0 downto 0);
        p_o_image1_8_7  : out    vl_logic_vector(1 downto 0);
        p_o_image1_8_1  : out    vl_logic_vector(1 downto 1);
        p_o_image1_8_2  : out    vl_logic_vector(1 downto 1);
        p_o_image1_8_3  : out    vl_logic_vector(1 downto 1);
        p_o_image1_8_4  : out    vl_logic_vector(1 downto 1);
        p_o_image1_8_5  : out    vl_logic_vector(1 downto 1);
        p_o_image1_8_6  : out    vl_logic_vector(1 downto 1);
        p_o_image1_7    : out    vl_logic_vector(2 downto 1);
        p_o_image1_1    : out    vl_logic_vector(2 downto 2);
        p_o_image1_2    : out    vl_logic_vector(2 downto 2);
        p_o_image1_3    : out    vl_logic_vector(2 downto 2);
        p_o_image1_4    : out    vl_logic_vector(2 downto 2);
        p_o_image1_5    : out    vl_logic_vector(2 downto 2);
        p_o_image1_6    : out    vl_logic_vector(2 downto 2);
        p_o_image2_9_7  : out    vl_logic_vector(1 downto 0);
        p_o_image2_9_1  : out    vl_logic_vector(0 downto 0);
        p_o_image2_9_2  : out    vl_logic_vector(0 downto 0);
        p_o_image2_9_3  : out    vl_logic_vector(0 downto 0);
        p_o_image2_9_4  : out    vl_logic_vector(0 downto 0);
        p_o_image2_9_5  : out    vl_logic_vector(0 downto 0);
        p_o_image2_9_6  : out    vl_logic_vector(0 downto 0);
        p_o_image2_8_7  : out    vl_logic_vector(1 downto 0);
        p_o_image2_8_1  : out    vl_logic_vector(1 downto 1);
        p_o_image2_8_2  : out    vl_logic_vector(1 downto 1);
        p_o_image2_8_3  : out    vl_logic_vector(1 downto 1);
        p_o_image2_8_4  : out    vl_logic_vector(1 downto 1);
        p_o_image2_8_5  : out    vl_logic_vector(1 downto 1);
        p_o_image2_8_6  : out    vl_logic_vector(1 downto 1);
        p_o_image2_7    : out    vl_logic_vector(2 downto 1);
        p_o_image2_1    : out    vl_logic_vector(2 downto 2);
        p_o_image2_2    : out    vl_logic_vector(2 downto 2);
        p_o_image2_3    : out    vl_logic_vector(2 downto 2);
        p_o_image2_4    : out    vl_logic_vector(2 downto 2);
        p_o_image2_5    : out    vl_logic_vector(2 downto 2);
        p_o_image2_6    : out    vl_logic_vector(2 downto 2);
        p_o_column      : out    vl_logic_vector(7 downto 0);
        p_debug_num_1   : out    vl_logic_vector(2 downto 0);
        p_o_mode        : out    vl_logic_vector(1 downto 0);
        p_debug_valid_modgen_and_1: in     vl_logic_vector(2 downto 2);
        p_i_valid_rtlc2_54_or_1: in     vl_logic_vector(2 downto 2);
        p_i_reset       : in     vl_logic;
        p_debug_num_0   : out    vl_logic_vector(2 downto 0);
        p_debug_num_2   : in     vl_logic_vector(7 downto 0);
        p_i_clock       : in     vl_logic;
        px1             : out    vl_logic;
        px23            : out    vl_logic;
        p_rtlc2n264     : out    vl_logic
    );
end memory_notri;
