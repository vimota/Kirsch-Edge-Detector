
library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.kirsch_utility_pkg.all;

entity kirsch is
	port(
		------------------------------------------
		-- main inputs and outputs
		i_clock    : in  std_logic;                      
		i_reset    : in  std_logic;                      
		i_valid    : in  std_logic;                 
		i_pixel    : in  std_logic_vector(7 downto 0);
		o_valid    : out std_logic;                 
		o_edge     : out std_logic;                      
		o_dir      : out std_logic_vector(2 downto 0);                      
		o_mode     : out std_logic_vector(1 downto 0);
		o_row      : out std_logic_vector(7 downto 0);
		o_column   : out std_logic_vector(7 downto 0);
		o_image0, o_image1, o_image2   : out image_type;
		------------------------------------------
		-- debugging inputs and outputs
		debug_key      : in  std_logic_vector( 3 downto 1) ; 
		debug_switch   : in  std_logic_vector(17 downto 0) ; 
		debug_led_red  : out std_logic_vector(17 downto 0) ; 
		debug_led_grn  : out std_logic_vector(5  downto 0) ; 
		debug_num_0    : out std_logic_vector(3 downto 0) ; 
		debug_num_1    : out std_logic_vector(3 downto 0) ; 
		debug_num_2    : out std_logic_vector(3 downto 0) ; 
		debug_num_3    : out std_logic_vector(3 downto 0) ; 
		debug_num_4    : out std_logic_vector(3 downto 0) ;
		debug_num_5    : out std_logic_vector(3 downto 0) 
		------------------------------------------
	);  
end entity;


architecture main of kirsch is
begin  
		-- instantiate memory
	u_memory : entity work.memory(main) port map 
	(
		i_valid  => i_valid,
		i_reset  => i_reset,
		i_pixel  => i_pixel,
		i_clock  => i_clock,
		-- o_valid  : out std_logic;
		-- o_mode   : out std_logic_vector(2 downto 0);
		o_column => o_column,
		o_image0 => o_image0,
		o_image1 => o_image1,
		o_image2 => o_image2,
		o_row    => o_row
	);


	debug_num_5 <= X"E";
	debug_num_4 <= X"C";
	debug_num_3 <= X"E";
	debug_num_2 <= X"3";
	debug_num_1 <= X"2";
	debug_num_0 <= X"7";

	debug_led_red <= (others => '0');
	debug_led_grn <= (others => '0');
	
end architecture;
