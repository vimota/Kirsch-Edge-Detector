//
// Verilog description for cell memory, 
// Mon Jul 21 14:16:47 2014
//
// Precision RTL Synthesis, 2008a.47//


module memory ( i_valid, i_reset, i_pixel, i_clock, o_valid, o_mode, o_column, 
                o_row, o_image0_0_, o_image0_1_, o_image0_2_, o_image1_0_, 
                o_image1_1_, o_image1_2_, o_image2_0_, o_image2_1_, o_image2_2_
                 ) ;

    input i_valid ;
    input i_reset ;
    input [7:0]i_pixel ;
    input i_clock ;
    output o_valid ;
    output [1:0]o_mode ;
    output [7:0]o_column ;
    output [7:0]o_row ;
    output [7:0]o_image0_0_ ;
    output [7:0]o_image0_1_ ;
    output [7:0]o_image0_2_ ;
    output [7:0]o_image1_0_ ;
    output [7:0]o_image1_1_ ;
    output [7:0]o_image1_2_ ;
    output [7:0]o_image2_0_ ;
    output [7:0]o_image2_1_ ;
    output [7:0]o_image2_2_ ;

    wire o_valid_dup0;
    wire [2:0]mem_wrn;
    wire [2:0]mem_wrn_current;
    wire first_bubble, busySignal, busySignalDelayed;
    wire [7:0]column;
    wire [7:0]row;
    wire [7:0]o_image1_dup0;
    wire o_image1_1__dup0_7_, o_image1_1__dup0_6_, o_image1_1__dup0_5_, 
         o_image1_1__dup0_4_, o_image1_1__dup0_3_, o_image1_1__dup0_2_, 
         o_image1_1__dup0_1_, o_image1_1__dup0_0_, o_image1_2__dup0_7_, 
         o_image1_2__dup0_6_, o_image1_2__dup0_5_, o_image1_2__dup0_4_, 
         o_image1_2__dup0_3_, o_image1_2__dup0_2_, o_image1_2__dup0_1_, 
         o_image1_2__dup0_0_;
    wire [7:0]o_image2_dup0;
    wire o_image2_1__dup0_7_, o_image2_1__dup0_6_, o_image2_1__dup0_5_, 
         o_image2_1__dup0_4_, o_image2_1__dup0_3_, o_image2_1__dup0_2_, 
         o_image2_1__dup0_1_, o_image2_1__dup0_0_, o_image2_2__dup0_7_, 
         o_image2_2__dup0_6_, o_image2_2__dup0_5_, o_image2_2__dup0_4_, 
         o_image2_2__dup0_3_, o_image2_2__dup0_2_, o_image2_2__dup0_1_, 
         o_image2_2__dup0_0_;
    wire [7:0]mem_q_0_;
    wire [7:0]mem_q_1_;
    wire [7:0]mem_q_2_;
    wire i_valid_int, i_reset_int;
    wire [7:0]i_pixel_int;
    wire i_clock_int;
    wire [1:0]o_mode_dup0;
    wire nx8852z1, nx15763z4, not_first_bubble, not_rtlc3_X_0_n252, nx47386z1, 
         nx15763z3, nx15763z2, nx16760z1;
    wire [7:0]buffer2_4n2ss1;
    wire nx60567z2, nx8852z2, nx33254z1, nx39109z3, nx41103z4, nx63578z4, 
         nx62359z4, nx8852z3, nx60567z1, nx5021z2, nx4024z2, nx3027z2, nx2030z2, 
         nx1033z2, nx36z2, nx64575z2, nx63578z2, nx55380z2, nx56377z2, nx57374z2, 
         nx58371z2, nx59368z2, nx60365z2, nx61362z2, nx62359z2, nx41103z1, 
         nx39109z2, nx8852z4, nx8852z6, nx8852z7, nx60567z3, nx60567z4, 
         nx60567z5, nx63578z3, nx62359z3, nx60567z6, nx41103z3, nx41103z2, 
         nx8852z5, nx57224z1, nx56227z1, nx55230z1, nx54233z1, nx53236z1, 
         nx52239z1, nx51242z1, nx50245z1, nx62359z1, nx61362z1, nx60365z1, 
         nx59368z1, nx58371z1, nx57374z1, nx56377z1, nx55380z1, nx63578z1, 
         nx64575z1, nx36z1, nx1033z1, nx2030z1, nx3027z1, nx4024z1, nx5021z1, 
         nx30938z1, nx31935z1, nx32932z1, nx33929z1, nx34926z1, nx35923z1, 
         nx36920z1, nx37917z1, nx36073z1, nx37070z1, nx38067z1, nx39064z1, 
         nx40061z1, nx41058z1, nx42055z1, nx43052z1, nx41208z1, nx42205z1, 
         nx43202z1, nx44199z1, nx45196z1, nx46193z1, nx47190z1, nx48187z1, 
         nx4207z1, nx3210z1, nx2213z1, nx1216z1, nx219z1, nx64758z1, nx63761z1, 
         nx62764z1, nx64608z1, nx63611z1, nx62614z1, nx61617z1, nx60620z1, 
         nx59623z1, nx58626z1, nx57629z1, nx59473z1, nx58476z1, nx57479z1, 
         nx56482z1, nx55485z1, nx54488z1, nx53491z1, nx52494z1, nx16335z1, 
         nx17332z1, nx18329z1, nx19326z1, nx20323z1, nx21320z1, nx22317z1, 
         nx23314z1, nx4657z1, nx5654z1, nx6651z1, nx7648z1, nx8645z1, nx9642z1, 
         nx10639z1, nx11636z1, nx39109z1, nx15763z1;
    wire [2386:0] xmplr_dummy ;




    modgen_counter_8_0 modgen_counter_row (.clock (i_clock_int), .q ({row[7],
                       row[6],row[5],row[4],row[3],row[2],row[1],row[0]}), .sclear (
                       nx8852z1), .cnt_en (not_rtlc3_X_0_n252), .p_rtlc6n55 (
                       nx8852z2), .p_i_reset_int (i_reset_int)) ;
    modgen_counter_8_1 modgen_counter_column (.clock (i_clock_int), .q ({
                       column[7],column[6],column[5],column[4],column[3],
                       column[2],column[1],column[0]}), .sclear (nx47386z1), .cnt_en (
                       first_bubble), .p_rtlc3n121 (nx8852z1), .p_i_valid_int (
                       i_valid_int)) ;
    ram_dq_8_0 u_mem1_mem (.wr_data1 ({i_pixel_int[7],i_pixel_int[6],
               i_pixel_int[5],i_pixel_int[4],i_pixel_int[3],i_pixel_int[2],
               i_pixel_int[1],i_pixel_int[0]}), .rd_data1 ({mem_q_0_[7],
               mem_q_0_[6],mem_q_0_[5],mem_q_0_[4],mem_q_0_[3],mem_q_0_[2],
               mem_q_0_[1],mem_q_0_[0]}), .addr1 ({column[7],column[6],column[5]
               ,column[4],column[3],column[2],column[1],column[0]}), .wr_clk1 (
               i_clock_int), .wr_ena1 (mem_wrn[0])) ;
    ram_dq_8_1 u_mem2_mem (.wr_data1 ({i_pixel_int[7],i_pixel_int[6],
               i_pixel_int[5],i_pixel_int[4],i_pixel_int[3],i_pixel_int[2],
               i_pixel_int[1],i_pixel_int[0]}), .rd_data1 ({mem_q_1_[7],
               mem_q_1_[6],mem_q_1_[5],mem_q_1_[4],mem_q_1_[3],mem_q_1_[2],
               mem_q_1_[1],mem_q_1_[0]}), .addr1 ({column[7],column[6],column[5]
               ,column[4],column[3],column[2],column[1],column[0]}), .wr_clk1 (
               i_clock_int), .wr_ena1 (mem_wrn[1])) ;
    ram_dq_8_2 u_mem3_mem (.wr_data1 ({i_pixel_int[7],i_pixel_int[6],
               i_pixel_int[5],i_pixel_int[4],i_pixel_int[3],i_pixel_int[2],
               i_pixel_int[1],i_pixel_int[0]}), .rd_data1 ({mem_q_2_[7],
               mem_q_2_[6],mem_q_2_[5],mem_q_2_[4],mem_q_2_[3],mem_q_2_[2],
               mem_q_2_[1],mem_q_2_[0]}), .addr1 ({column[7],column[6],column[5]
               ,column[4],column[3],column[2],column[1],column[0]}), .wr_clk1 (
               i_clock_int), .wr_ena1 (mem_wrn[2])) ;
    assign o_mode_dup0[1] = ~i_reset_int ;
    assign not_first_bubble = ~first_bubble ;
    cycloneii_lcell_ff reg_out_o_row_obuf_7_ (.regout (nx23314z1), .datain (
                       row[7]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_row_obuf_6_ (.regout (nx22317z1), .datain (
                       row[6]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_row_obuf_5_ (.regout (nx21320z1), .datain (
                       row[5]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_row_obuf_4_ (.regout (nx20323z1), .datain (
                       row[4]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_row_obuf_3_ (.regout (nx19326z1), .datain (
                       row[3]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_row_obuf_2_ (.regout (nx18329z1), .datain (
                       row[2]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_row_obuf_1_ (.regout (nx17332z1), .datain (
                       row[1]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_row_obuf_0_ (.regout (nx16335z1), .datain (
                       row[0]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), 
                       .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__7_ (.regout (nx37917z1), .datain (
                       o_image2_2__dup0_7_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__6_ (.regout (nx36920z1), .datain (
                       o_image2_2__dup0_6_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__5_ (.regout (nx35923z1), .datain (
                       o_image2_2__dup0_5_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__4_ (.regout (nx34926z1), .datain (
                       o_image2_2__dup0_4_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__3_ (.regout (nx33929z1), .datain (
                       o_image2_2__dup0_3_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__2_ (.regout (nx32932z1), .datain (
                       o_image2_2__dup0_2_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__1_ (.regout (nx31935z1), .datain (
                       o_image2_2__dup0_1_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_2__0_ (.regout (nx30938z1), .datain (
                       o_image2_2__dup0_0_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__7_ (.regout (nx43052z1), .datain (
                       o_image2_1__dup0_7_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__6_ (.regout (nx42055z1), .datain (
                       o_image2_1__dup0_6_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__5_ (.regout (nx41058z1), .datain (
                       o_image2_1__dup0_5_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__4_ (.regout (nx40061z1), .datain (
                       o_image2_1__dup0_4_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__3_ (.regout (nx39064z1), .datain (
                       o_image2_1__dup0_3_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__2_ (.regout (nx38067z1), .datain (
                       o_image2_1__dup0_2_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__1_ (.regout (nx37070z1), .datain (
                       o_image2_1__dup0_1_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_1__0_ (.regout (nx36073z1), .datain (
                       o_image2_1__dup0_0_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__7_ (.regout (nx48187z1), .datain (
                       o_image2_dup0[7]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__6_ (.regout (nx47190z1), .datain (
                       o_image2_dup0[6]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__5_ (.regout (nx46193z1), .datain (
                       o_image2_dup0[5]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__4_ (.regout (nx45196z1), .datain (
                       o_image2_dup0[4]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__3_ (.regout (nx44199z1), .datain (
                       o_image2_dup0[3]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__2_ (.regout (nx43202z1), .datain (
                       o_image2_dup0[2]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__1_ (.regout (nx42205z1), .datain (
                       o_image2_dup0[1]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image1_obuf_0__0_ (.regout (nx41208z1), .datain (
                       o_image2_dup0[0]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__7_ (.regout (nx62764z1), .datain (
                       o_image1_2__dup0_7_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__6_ (.regout (nx63761z1), .datain (
                       o_image1_2__dup0_6_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__5_ (.regout (nx64758z1), .datain (
                       o_image1_2__dup0_5_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__4_ (.regout (nx219z1), .datain (
                       o_image1_2__dup0_4_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__3_ (.regout (nx1216z1), .datain (
                       o_image1_2__dup0_3_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__2_ (.regout (nx2213z1), .datain (
                       o_image1_2__dup0_2_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__1_ (.regout (nx3210z1), .datain (
                       o_image1_2__dup0_1_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_2__0_ (.regout (nx4207z1), .datain (
                       o_image1_2__dup0_0_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__7_ (.regout (nx57629z1), .datain (
                       o_image1_1__dup0_7_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__6_ (.regout (nx58626z1), .datain (
                       o_image1_1__dup0_6_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__5_ (.regout (nx59623z1), .datain (
                       o_image1_1__dup0_5_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__4_ (.regout (nx60620z1), .datain (
                       o_image1_1__dup0_4_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__3_ (.regout (nx61617z1), .datain (
                       o_image1_1__dup0_3_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__2_ (.regout (nx62614z1), .datain (
                       o_image1_1__dup0_2_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__1_ (.regout (nx63611z1), .datain (
                       o_image1_1__dup0_1_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_1__0_ (.regout (nx64608z1), .datain (
                       o_image1_1__dup0_0_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__7_ (.regout (nx52494z1), .datain (
                       o_image1_dup0[7]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__6_ (.regout (nx53491z1), .datain (
                       o_image1_dup0[6]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__5_ (.regout (nx54488z1), .datain (
                       o_image1_dup0[5]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__4_ (.regout (nx55485z1), .datain (
                       o_image1_dup0[4]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__3_ (.regout (nx56482z1), .datain (
                       o_image1_dup0[3]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__2_ (.regout (nx57479z1), .datain (
                       o_image1_dup0[2]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__1_ (.regout (nx58476z1), .datain (
                       o_image1_dup0[1]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_image0_obuf_0__0_ (.regout (nx59473z1), .datain (
                       o_image1_dup0[0]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_7_ (.regout (nx11636z1), .datain (
                       column[7]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_6_ (.regout (nx10639z1), .datain (
                       column[6]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_5_ (.regout (nx9642z1), .datain (
                       column[5]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_4_ (.regout (nx8645z1), .datain (
                       column[4]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_3_ (.regout (nx7648z1), .datain (
                       column[3]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_2_ (.regout (nx6651z1), .datain (
                       column[2]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_1_ (.regout (nx5654z1), .datain (
                       column[1]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_out_o_column_obuf_0_ (.regout (nx4657z1), .datain (
                       column[0]), .sdata (1'b0), .clk (i_clock_int), .ena (1'b1
                       ), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_o_valid (.regout (o_valid_dup0), .datain (nx60567z1)
                       , .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), .aclr (
                       1'b0), .sclr (not_first_bubble), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_mem_wrn_current_2_ (.regout (mem_wrn_current[2]), .datain (
                       mem_wrn_current[1]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       nx41103z1), .aclr (1'b0), .sclr (nx41103z4), .sload (1'b0
                       )) ;
    cycloneii_lcell_ff reg_mem_wrn_current_1_ (.regout (mem_wrn_current[1]), .datain (
                       mem_wrn_current[0]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       nx41103z1), .aclr (1'b0), .sclr (nx41103z4), .sload (1'b0
                       )) ;
    assign nx39109z1 = 1 ;
    cycloneii_lcell_ff reg_mem_wrn_current_0_ (.regout (mem_wrn_current[0]), .datain (
                       mem_wrn_current[2]), .sdata (nx39109z1), .clk (
                       i_clock_int), .ena (nx39109z2), .aclr (1'b0), .sclr (
                       nx8852z1), .sload (nx39109z3)) ;
    cycloneii_lcell_ff reg_mem_wrn_2_ (.regout (mem_wrn[2]), .datain (
                       mem_wrn_current[2]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       1'b1), .aclr (1'b0), .sclr (nx16760z1), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_mem_wrn_1_ (.regout (mem_wrn[1]), .datain (
                       mem_wrn_current[1]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       1'b1), .aclr (1'b0), .sclr (nx16760z1), .sload (1'b0)) ;
    assign nx15763z1 = 1 ;
    cycloneii_lcell_ff reg_mem_wrn_0_ (.regout (mem_wrn[0]), .datain (
                       mem_wrn_current[0]), .sdata (nx15763z1), .clk (
                       i_clock_int), .ena (1'b1), .aclr (1'b0), .sclr (nx15763z2
                       ), .sload (nx15763z3)) ;
    cycloneii_lcell_ff reg_in_i_valid_ibuf (.regout (first_bubble), .datain (
                       i_valid_int), .sdata (1'b0), .clk (i_clock_int), .ena (
                       1'b1), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_busySignalDelayed (.regout (busySignalDelayed), .datain (
                       busySignal), .sdata (1'b0), .clk (i_clock_int), .ena (
                       1'b1), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_busySignal (.regout (busySignal), .datain (nx33254z1)
                       , .sdata (1'b0), .clk (i_clock_int), .ena (1'b1), .aclr (
                       1'b0), .sclr (nx8852z2), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_buffer2_2__7_ (.regout (o_image2_2__dup0_7_), .datain (
                       nx57224z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_2__6_ (.regout (o_image2_2__dup0_6_), .datain (
                       nx56227z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_2__5_ (.regout (o_image2_2__dup0_5_), .datain (
                       nx55230z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_2__4_ (.regout (o_image2_2__dup0_4_), .datain (
                       nx54233z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_2__3_ (.regout (o_image2_2__dup0_3_), .datain (
                       nx53236z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_2__2_ (.regout (o_image2_2__dup0_2_), .datain (
                       nx52239z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_2__1_ (.regout (o_image2_2__dup0_1_), .datain (
                       nx51242z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_2__0_ (.regout (o_image2_2__dup0_0_), .datain (
                       nx50245z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__7_ (.regout (o_image2_1__dup0_7_), .datain (
                       nx62359z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__6_ (.regout (o_image2_1__dup0_6_), .datain (
                       nx61362z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__5_ (.regout (o_image2_1__dup0_5_), .datain (
                       nx60365z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__4_ (.regout (o_image2_1__dup0_4_), .datain (
                       nx59368z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__3_ (.regout (o_image2_1__dup0_3_), .datain (
                       nx58371z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__2_ (.regout (o_image2_1__dup0_2_), .datain (
                       nx57374z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__1_ (.regout (o_image2_1__dup0_1_), .datain (
                       nx56377z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_1__0_ (.regout (o_image2_1__dup0_0_), .datain (
                       nx55380z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__7_ (.regout (o_image2_dup0[7]), .datain (
                       nx63578z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__6_ (.regout (o_image2_dup0[6]), .datain (
                       nx64575z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__5_ (.regout (o_image2_dup0[5]), .datain (
                       nx36z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__4_ (.regout (o_image2_dup0[4]), .datain (
                       nx1033z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__3_ (.regout (o_image2_dup0[3]), .datain (
                       nx2030z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__2_ (.regout (o_image2_dup0[2]), .datain (
                       nx3027z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__1_ (.regout (o_image2_dup0[1]), .datain (
                       nx4024z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer2_0__0_ (.regout (o_image2_dup0[0]), .datain (
                       nx5021z1), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_2__7_ (.regout (o_image1_2__dup0_7_), .datain (
                       o_image2_2__dup0_7_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_2__6_ (.regout (o_image1_2__dup0_6_), .datain (
                       o_image2_2__dup0_6_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_2__5_ (.regout (o_image1_2__dup0_5_), .datain (
                       o_image2_2__dup0_5_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_2__4_ (.regout (o_image1_2__dup0_4_), .datain (
                       o_image2_2__dup0_4_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_2__3_ (.regout (o_image1_2__dup0_3_), .datain (
                       o_image2_2__dup0_3_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_2__2_ (.regout (o_image1_2__dup0_2_), .datain (
                       o_image2_2__dup0_2_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_2__1_ (.regout (o_image1_2__dup0_1_), .datain (
                       o_image2_2__dup0_1_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_2__0_ (.regout (o_image1_2__dup0_0_), .datain (
                       o_image2_2__dup0_0_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__7_ (.regout (o_image1_1__dup0_7_), .datain (
                       o_image2_1__dup0_7_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__6_ (.regout (o_image1_1__dup0_6_), .datain (
                       o_image2_1__dup0_6_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__5_ (.regout (o_image1_1__dup0_5_), .datain (
                       o_image2_1__dup0_5_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__4_ (.regout (o_image1_1__dup0_4_), .datain (
                       o_image2_1__dup0_4_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__3_ (.regout (o_image1_1__dup0_3_), .datain (
                       o_image2_1__dup0_3_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__2_ (.regout (o_image1_1__dup0_2_), .datain (
                       o_image2_1__dup0_2_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__1_ (.regout (o_image1_1__dup0_1_), .datain (
                       o_image2_1__dup0_1_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_1__0_ (.regout (o_image1_1__dup0_0_), .datain (
                       o_image2_1__dup0_0_), .sdata (1'b0), .clk (i_clock_int), 
                       .ena (first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (
                       1'b0)) ;
    cycloneii_lcell_ff reg_buffer1_0__7_ (.regout (o_image1_dup0[7]), .datain (
                       o_image2_dup0[7]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_0__6_ (.regout (o_image1_dup0[6]), .datain (
                       o_image2_dup0[6]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_0__5_ (.regout (o_image1_dup0[5]), .datain (
                       o_image2_dup0[5]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_0__4_ (.regout (o_image1_dup0[4]), .datain (
                       o_image2_dup0[4]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_0__3_ (.regout (o_image1_dup0[3]), .datain (
                       o_image2_dup0[3]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_0__2_ (.regout (o_image1_dup0[2]), .datain (
                       o_image2_dup0[2]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_0__1_ (.regout (o_image1_dup0[1]), .datain (
                       o_image2_dup0[1]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_lcell_ff reg_buffer1_0__0_ (.regout (o_image1_dup0[0]), .datain (
                       o_image2_dup0[0]), .sdata (1'b0), .clk (i_clock_int), .ena (
                       first_bubble), .aclr (1'b0), .sclr (1'b0), .sload (1'b0)
                       ) ;
    cycloneii_io o_valid_obuf (.padio (o_valid), .datain (o_valid_dup0), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam o_valid_obuf.operation_mode = "output";
                 
                 defparam o_valid_obuf.output_register_mode = "none";
                 
                 defparam o_valid_obuf.tie_off_output_clock_enable = "false";
                 
                 defparam o_valid_obuf.oe_register_mode = "none";
                 
                 defparam o_valid_obuf.tie_off_oe_clock_enable = "false";
                 
                 defparam o_valid_obuf.input_register_mode = "none";
    cycloneii_io o_mode_obuf_1_ (.padio (o_mode[1]), .datain (o_mode_dup0[1]), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam o_mode_obuf_1_.operation_mode = "output";
                 
                 defparam o_mode_obuf_1_.output_register_mode = "none";
                 
                 defparam o_mode_obuf_1_.tie_off_output_clock_enable = "false";
                 
                 defparam o_mode_obuf_1_.oe_register_mode = "none";
                 
                 defparam o_mode_obuf_1_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_mode_obuf_1_.input_register_mode = "none";
    cycloneii_io o_mode_obuf_0_ (.padio (o_mode[0]), .datain (o_mode_dup0[0]), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam o_mode_obuf_0_.operation_mode = "output";
                 
                 defparam o_mode_obuf_0_.output_register_mode = "none";
                 
                 defparam o_mode_obuf_0_.tie_off_output_clock_enable = "false";
                 
                 defparam o_mode_obuf_0_.oe_register_mode = "none";
                 
                 defparam o_mode_obuf_0_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_mode_obuf_0_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__7_ (.padio (o_image2_2_[7]), .datain (
                 o_image2_2__dup0_7_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__7_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__7_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__7_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__7_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__7_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__7_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__6_ (.padio (o_image2_2_[6]), .datain (
                 o_image2_2__dup0_6_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__6_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__6_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__6_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__6_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__6_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__6_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__5_ (.padio (o_image2_2_[5]), .datain (
                 o_image2_2__dup0_5_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__5_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__5_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__5_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__5_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__5_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__5_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__4_ (.padio (o_image2_2_[4]), .datain (
                 o_image2_2__dup0_4_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__4_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__4_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__4_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__4_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__4_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__4_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__3_ (.padio (o_image2_2_[3]), .datain (
                 o_image2_2__dup0_3_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__3_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__3_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__3_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__3_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__3_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__3_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__2_ (.padio (o_image2_2_[2]), .datain (
                 o_image2_2__dup0_2_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__2_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__2_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__2_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__2_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__2_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__2_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__1_ (.padio (o_image2_2_[1]), .datain (
                 o_image2_2__dup0_1_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__1_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__1_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__1_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__1_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__1_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__1_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_2__0_ (.padio (o_image2_2_[0]), .datain (
                 o_image2_2__dup0_0_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_2__0_.operation_mode = "output";
                 
                 defparam o_image2_obuf_2__0_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_2__0_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__0_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_2__0_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_2__0_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__7_ (.padio (o_image2_1_[7]), .datain (
                 o_image2_1__dup0_7_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__7_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__7_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__7_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__7_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__7_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__7_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__6_ (.padio (o_image2_1_[6]), .datain (
                 o_image2_1__dup0_6_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__6_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__6_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__6_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__6_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__6_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__6_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__5_ (.padio (o_image2_1_[5]), .datain (
                 o_image2_1__dup0_5_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__5_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__5_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__5_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__5_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__5_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__5_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__4_ (.padio (o_image2_1_[4]), .datain (
                 o_image2_1__dup0_4_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__4_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__4_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__4_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__4_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__4_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__4_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__3_ (.padio (o_image2_1_[3]), .datain (
                 o_image2_1__dup0_3_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__3_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__3_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__3_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__3_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__3_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__3_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__2_ (.padio (o_image2_1_[2]), .datain (
                 o_image2_1__dup0_2_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__2_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__2_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__2_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__2_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__2_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__2_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__1_ (.padio (o_image2_1_[1]), .datain (
                 o_image2_1__dup0_1_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__1_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__1_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__1_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__1_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__1_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__1_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_1__0_ (.padio (o_image2_1_[0]), .datain (
                 o_image2_1__dup0_0_), .oe (1'b1), .outclk (1'b0), .outclkena (
                 1'b1), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_1__0_.operation_mode = "output";
                 
                 defparam o_image2_obuf_1__0_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_1__0_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__0_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_1__0_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_1__0_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__7_ (.padio (o_image2_0_[7]), .datain (
                 o_image2_dup0[7]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__7_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__7_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__7_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__7_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__7_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__7_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__6_ (.padio (o_image2_0_[6]), .datain (
                 o_image2_dup0[6]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__6_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__6_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__6_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__6_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__6_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__6_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__5_ (.padio (o_image2_0_[5]), .datain (
                 o_image2_dup0[5]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__5_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__5_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__5_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__5_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__5_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__5_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__4_ (.padio (o_image2_0_[4]), .datain (
                 o_image2_dup0[4]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__4_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__4_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__4_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__4_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__4_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__4_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__3_ (.padio (o_image2_0_[3]), .datain (
                 o_image2_dup0[3]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__3_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__3_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__3_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__3_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__3_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__3_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__2_ (.padio (o_image2_0_[2]), .datain (
                 o_image2_dup0[2]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__2_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__2_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__2_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__2_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__2_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__2_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__1_ (.padio (o_image2_0_[1]), .datain (
                 o_image2_dup0[1]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__1_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__1_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__1_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__1_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__1_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__1_.input_register_mode = "none";
    cycloneii_io o_image2_obuf_0__0_ (.padio (o_image2_0_[0]), .datain (
                 o_image2_dup0[0]), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1
                 ), .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 
                 defparam o_image2_obuf_0__0_.operation_mode = "output";
                 
                 defparam o_image2_obuf_0__0_.output_register_mode = "none";
                 
                 defparam o_image2_obuf_0__0_.tie_off_output_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__0_.oe_register_mode = "none";
                 
                 defparam o_image2_obuf_0__0_.tie_off_oe_clock_enable = "false";
                 
                 defparam o_image2_obuf_0__0_.input_register_mode = "none";
    cycloneii_io ix13876z43919 (.combout (i_valid_int), .padio (i_valid), .datain (
                 1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (
                 1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix13876z43919.operation_mode = "input";
                 
                 defparam ix13876z43919.output_register_mode = "none";
                 
                 defparam ix13876z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix13876z43919.oe_register_mode = "none";
                 
                 defparam ix13876z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix13876z43919.input_register_mode = "none";
    cycloneii_io ix11636z43919 (.padio (o_column[7]), .datain (nx11636z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix11636z43919.operation_mode = "output";
                 
                 defparam ix11636z43919.output_register_mode = "none";
                 
                 defparam ix11636z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix11636z43919.oe_register_mode = "none";
                 
                 defparam ix11636z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix11636z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix5021z52923 (.combout (nx5021z1), .dataa (1'b1), .datab (
                         nx5021z2), .datac (mem_q_0_[0]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix5021z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix10639z43919 (.padio (o_column[6]), .datain (nx10639z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix10639z43919.operation_mode = "output";
                 
                 defparam ix10639z43919.output_register_mode = "none";
                 
                 defparam ix10639z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix10639z43919.oe_register_mode = "none";
                 
                 defparam ix10639z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix10639z43919.input_register_mode = "none";
    cycloneii_io ix9642z43919 (.padio (o_column[5]), .datain (nx9642z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix9642z43919.operation_mode = "output";
                 
                 defparam ix9642z43919.output_register_mode = "none";
                 
                 defparam ix9642z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix9642z43919.oe_register_mode = "none";
                 
                 defparam ix9642z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix9642z43919.input_register_mode = "none";
    cycloneii_io ix8645z43919 (.padio (o_column[4]), .datain (nx8645z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix8645z43919.operation_mode = "output";
                 
                 defparam ix8645z43919.output_register_mode = "none";
                 
                 defparam ix8645z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix8645z43919.oe_register_mode = "none";
                 
                 defparam ix8645z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix8645z43919.input_register_mode = "none";
    cycloneii_io ix7648z43919 (.padio (o_column[3]), .datain (nx7648z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix7648z43919.operation_mode = "output";
                 
                 defparam ix7648z43919.output_register_mode = "none";
                 
                 defparam ix7648z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix7648z43919.oe_register_mode = "none";
                 
                 defparam ix7648z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix7648z43919.input_register_mode = "none";
    cycloneii_io ix6651z43919 (.padio (o_column[2]), .datain (nx6651z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix6651z43919.operation_mode = "output";
                 
                 defparam ix6651z43919.output_register_mode = "none";
                 
                 defparam ix6651z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix6651z43919.oe_register_mode = "none";
                 
                 defparam ix6651z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix6651z43919.input_register_mode = "none";
    cycloneii_io ix5654z43919 (.padio (o_column[1]), .datain (nx5654z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix5654z43919.operation_mode = "output";
                 
                 defparam ix5654z43919.output_register_mode = "none";
                 
                 defparam ix5654z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix5654z43919.oe_register_mode = "none";
                 
                 defparam ix5654z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix5654z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix4024z52923 (.combout (nx4024z1), .dataa (1'b1), .datab (
                         nx4024z2), .datac (mem_q_0_[1]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix4024z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix4657z43919 (.padio (o_column[0]), .datain (nx4657z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix4657z43919.operation_mode = "output";
                 
                 defparam ix4657z43919.output_register_mode = "none";
                 
                 defparam ix4657z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix4657z43919.oe_register_mode = "none";
                 
                 defparam ix4657z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix4657z43919.input_register_mode = "none";
    cycloneii_io ix23314z43919 (.padio (o_row[7]), .datain (nx23314z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix23314z43919.operation_mode = "output";
                 
                 defparam ix23314z43919.output_register_mode = "none";
                 
                 defparam ix23314z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix23314z43919.oe_register_mode = "none";
                 
                 defparam ix23314z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix23314z43919.input_register_mode = "none";
    cycloneii_io ix22317z43919 (.padio (o_row[6]), .datain (nx22317z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix22317z43919.operation_mode = "output";
                 
                 defparam ix22317z43919.output_register_mode = "none";
                 
                 defparam ix22317z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix22317z43919.oe_register_mode = "none";
                 
                 defparam ix22317z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix22317z43919.input_register_mode = "none";
    cycloneii_io ix21320z43919 (.padio (o_row[5]), .datain (nx21320z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix21320z43919.operation_mode = "output";
                 
                 defparam ix21320z43919.output_register_mode = "none";
                 
                 defparam ix21320z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix21320z43919.oe_register_mode = "none";
                 
                 defparam ix21320z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix21320z43919.input_register_mode = "none";
    cycloneii_io ix20323z43919 (.padio (o_row[4]), .datain (nx20323z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix20323z43919.operation_mode = "output";
                 
                 defparam ix20323z43919.output_register_mode = "none";
                 
                 defparam ix20323z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix20323z43919.oe_register_mode = "none";
                 
                 defparam ix20323z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix20323z43919.input_register_mode = "none";
    cycloneii_io ix19326z43919 (.padio (o_row[3]), .datain (nx19326z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix19326z43919.operation_mode = "output";
                 
                 defparam ix19326z43919.output_register_mode = "none";
                 
                 defparam ix19326z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix19326z43919.oe_register_mode = "none";
                 
                 defparam ix19326z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix19326z43919.input_register_mode = "none";
    cycloneii_io ix18329z43919 (.padio (o_row[2]), .datain (nx18329z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix18329z43919.operation_mode = "output";
                 
                 defparam ix18329z43919.output_register_mode = "none";
                 
                 defparam ix18329z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix18329z43919.oe_register_mode = "none";
                 
                 defparam ix18329z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix18329z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix3027z52923 (.combout (nx3027z1), .dataa (1'b1), .datab (
                         nx3027z2), .datac (mem_q_0_[2]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix3027z52923.lut_mask = 16'hf0cc;
    cycloneii_lcell_comb ix2030z52923 (.combout (nx2030z1), .dataa (1'b1), .datab (
                         nx2030z2), .datac (mem_q_0_[3]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix2030z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix17332z43919 (.padio (o_row[1]), .datain (nx17332z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix17332z43919.operation_mode = "output";
                 
                 defparam ix17332z43919.output_register_mode = "none";
                 
                 defparam ix17332z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix17332z43919.oe_register_mode = "none";
                 
                 defparam ix17332z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix17332z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix1033z52923 (.combout (nx1033z1), .dataa (1'b1), .datab (
                         nx1033z2), .datac (mem_q_0_[4]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix1033z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix16335z43919 (.padio (o_row[0]), .datain (nx16335z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix16335z43919.operation_mode = "output";
                 
                 defparam ix16335z43919.output_register_mode = "none";
                 
                 defparam ix16335z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix16335z43919.oe_register_mode = "none";
                 
                 defparam ix16335z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix16335z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix36z52923 (.combout (nx36z1), .dataa (1'b1), .datab (
                         nx36z2), .datac (mem_q_0_[5]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix36z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix52494z43919 (.padio (o_image0_0_[7]), .datain (nx52494z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix52494z43919.operation_mode = "output";
                 
                 defparam ix52494z43919.output_register_mode = "none";
                 
                 defparam ix52494z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix52494z43919.oe_register_mode = "none";
                 
                 defparam ix52494z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix52494z43919.input_register_mode = "none";
    cycloneii_io ix53491z43919 (.padio (o_image0_0_[6]), .datain (nx53491z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix53491z43919.operation_mode = "output";
                 
                 defparam ix53491z43919.output_register_mode = "none";
                 
                 defparam ix53491z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix53491z43919.oe_register_mode = "none";
                 
                 defparam ix53491z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix53491z43919.input_register_mode = "none";
    cycloneii_io ix54488z43919 (.padio (o_image0_0_[5]), .datain (nx54488z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix54488z43919.operation_mode = "output";
                 
                 defparam ix54488z43919.output_register_mode = "none";
                 
                 defparam ix54488z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix54488z43919.oe_register_mode = "none";
                 
                 defparam ix54488z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix54488z43919.input_register_mode = "none";
    cycloneii_io ix55485z43919 (.padio (o_image0_0_[4]), .datain (nx55485z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix55485z43919.operation_mode = "output";
                 
                 defparam ix55485z43919.output_register_mode = "none";
                 
                 defparam ix55485z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix55485z43919.oe_register_mode = "none";
                 
                 defparam ix55485z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix55485z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix64575z52923 (.combout (nx64575z1), .dataa (1'b1), .datab (
                         nx64575z2), .datac (mem_q_0_[6]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix64575z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix56482z43919 (.padio (o_image0_0_[3]), .datain (nx56482z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix56482z43919.operation_mode = "output";
                 
                 defparam ix56482z43919.output_register_mode = "none";
                 
                 defparam ix56482z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix56482z43919.oe_register_mode = "none";
                 
                 defparam ix56482z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix56482z43919.input_register_mode = "none";
    cycloneii_io ix57479z43919 (.padio (o_image0_0_[2]), .datain (nx57479z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix57479z43919.operation_mode = "output";
                 
                 defparam ix57479z43919.output_register_mode = "none";
                 
                 defparam ix57479z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix57479z43919.oe_register_mode = "none";
                 
                 defparam ix57479z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix57479z43919.input_register_mode = "none";
    cycloneii_io ix58476z43919 (.padio (o_image0_0_[1]), .datain (nx58476z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix58476z43919.operation_mode = "output";
                 
                 defparam ix58476z43919.output_register_mode = "none";
                 
                 defparam ix58476z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix58476z43919.oe_register_mode = "none";
                 
                 defparam ix58476z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix58476z43919.input_register_mode = "none";
    cycloneii_io ix59473z43919 (.padio (o_image0_0_[0]), .datain (nx59473z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix59473z43919.operation_mode = "output";
                 
                 defparam ix59473z43919.output_register_mode = "none";
                 
                 defparam ix59473z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix59473z43919.oe_register_mode = "none";
                 
                 defparam ix59473z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix59473z43919.input_register_mode = "none";
    cycloneii_io ix57629z43919 (.padio (o_image0_1_[7]), .datain (nx57629z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix57629z43919.operation_mode = "output";
                 
                 defparam ix57629z43919.output_register_mode = "none";
                 
                 defparam ix57629z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix57629z43919.oe_register_mode = "none";
                 
                 defparam ix57629z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix57629z43919.input_register_mode = "none";
    cycloneii_io ix58626z43919 (.padio (o_image0_1_[6]), .datain (nx58626z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix58626z43919.operation_mode = "output";
                 
                 defparam ix58626z43919.output_register_mode = "none";
                 
                 defparam ix58626z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix58626z43919.oe_register_mode = "none";
                 
                 defparam ix58626z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix58626z43919.input_register_mode = "none";
    cycloneii_io ix59623z43919 (.padio (o_image0_1_[5]), .datain (nx59623z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix59623z43919.operation_mode = "output";
                 
                 defparam ix59623z43919.output_register_mode = "none";
                 
                 defparam ix59623z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix59623z43919.oe_register_mode = "none";
                 
                 defparam ix59623z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix59623z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix63578z52923 (.combout (nx63578z1), .dataa (1'b1), .datab (
                         nx63578z2), .datac (mem_q_0_[7]), .datad (nx63578z4), .cin (
                         1'b0)) ;
                         defparam ix63578z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix60620z43919 (.padio (o_image0_1_[4]), .datain (nx60620z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix60620z43919.operation_mode = "output";
                 
                 defparam ix60620z43919.output_register_mode = "none";
                 
                 defparam ix60620z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix60620z43919.oe_register_mode = "none";
                 
                 defparam ix60620z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix60620z43919.input_register_mode = "none";
    cycloneii_io ix61617z43919 (.padio (o_image0_1_[3]), .datain (nx61617z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix61617z43919.operation_mode = "output";
                 
                 defparam ix61617z43919.output_register_mode = "none";
                 
                 defparam ix61617z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix61617z43919.oe_register_mode = "none";
                 
                 defparam ix61617z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix61617z43919.input_register_mode = "none";
    cycloneii_io ix62614z43919 (.padio (o_image0_1_[2]), .datain (nx62614z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix62614z43919.operation_mode = "output";
                 
                 defparam ix62614z43919.output_register_mode = "none";
                 
                 defparam ix62614z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix62614z43919.oe_register_mode = "none";
                 
                 defparam ix62614z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix62614z43919.input_register_mode = "none";
    cycloneii_io ix63611z43919 (.padio (o_image0_1_[1]), .datain (nx63611z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix63611z43919.operation_mode = "output";
                 
                 defparam ix63611z43919.output_register_mode = "none";
                 
                 defparam ix63611z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix63611z43919.oe_register_mode = "none";
                 
                 defparam ix63611z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix63611z43919.input_register_mode = "none";
    cycloneii_io ix64608z43919 (.padio (o_image0_1_[0]), .datain (nx64608z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix64608z43919.operation_mode = "output";
                 
                 defparam ix64608z43919.output_register_mode = "none";
                 
                 defparam ix64608z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix64608z43919.oe_register_mode = "none";
                 
                 defparam ix64608z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix64608z43919.input_register_mode = "none";
    cycloneii_io ix62764z43919 (.padio (o_image0_2_[7]), .datain (nx62764z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix62764z43919.operation_mode = "output";
                 
                 defparam ix62764z43919.output_register_mode = "none";
                 
                 defparam ix62764z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix62764z43919.oe_register_mode = "none";
                 
                 defparam ix62764z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix62764z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix55380z52923 (.combout (nx55380z1), .dataa (1'b1), .datab (
                         nx55380z2), .datac (mem_q_1_[0]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix55380z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix63761z43919 (.padio (o_image0_2_[6]), .datain (nx63761z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix63761z43919.operation_mode = "output";
                 
                 defparam ix63761z43919.output_register_mode = "none";
                 
                 defparam ix63761z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix63761z43919.oe_register_mode = "none";
                 
                 defparam ix63761z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix63761z43919.input_register_mode = "none";
    cycloneii_io ix64758z43919 (.padio (o_image0_2_[5]), .datain (nx64758z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix64758z43919.operation_mode = "output";
                 
                 defparam ix64758z43919.output_register_mode = "none";
                 
                 defparam ix64758z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix64758z43919.oe_register_mode = "none";
                 
                 defparam ix64758z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix64758z43919.input_register_mode = "none";
    cycloneii_io ix219z43919 (.padio (o_image0_2_[4]), .datain (nx219z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix219z43919.operation_mode = "output";
                 
                 defparam ix219z43919.output_register_mode = "none";
                 
                 defparam ix219z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix219z43919.oe_register_mode = "none";
                 
                 defparam ix219z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix219z43919.input_register_mode = "none";
    cycloneii_io ix1216z43919 (.padio (o_image0_2_[3]), .datain (nx1216z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix1216z43919.operation_mode = "output";
                 
                 defparam ix1216z43919.output_register_mode = "none";
                 
                 defparam ix1216z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix1216z43919.oe_register_mode = "none";
                 
                 defparam ix1216z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix1216z43919.input_register_mode = "none";
    cycloneii_io ix2213z43919 (.padio (o_image0_2_[2]), .datain (nx2213z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix2213z43919.operation_mode = "output";
                 
                 defparam ix2213z43919.output_register_mode = "none";
                 
                 defparam ix2213z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix2213z43919.oe_register_mode = "none";
                 
                 defparam ix2213z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix2213z43919.input_register_mode = "none";
    cycloneii_io ix3210z43919 (.padio (o_image0_2_[1]), .datain (nx3210z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix3210z43919.operation_mode = "output";
                 
                 defparam ix3210z43919.output_register_mode = "none";
                 
                 defparam ix3210z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix3210z43919.oe_register_mode = "none";
                 
                 defparam ix3210z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix3210z43919.input_register_mode = "none";
    cycloneii_io ix4207z43919 (.padio (o_image0_2_[0]), .datain (nx4207z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix4207z43919.operation_mode = "output";
                 
                 defparam ix4207z43919.output_register_mode = "none";
                 
                 defparam ix4207z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix4207z43919.oe_register_mode = "none";
                 
                 defparam ix4207z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix4207z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix56377z52923 (.combout (nx56377z1), .dataa (1'b1), .datab (
                         nx56377z2), .datac (mem_q_1_[1]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix56377z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix48187z43919 (.padio (o_image1_0_[7]), .datain (nx48187z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix48187z43919.operation_mode = "output";
                 
                 defparam ix48187z43919.output_register_mode = "none";
                 
                 defparam ix48187z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix48187z43919.oe_register_mode = "none";
                 
                 defparam ix48187z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix48187z43919.input_register_mode = "none";
    cycloneii_io ix47190z43919 (.padio (o_image1_0_[6]), .datain (nx47190z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix47190z43919.operation_mode = "output";
                 
                 defparam ix47190z43919.output_register_mode = "none";
                 
                 defparam ix47190z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix47190z43919.oe_register_mode = "none";
                 
                 defparam ix47190z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix47190z43919.input_register_mode = "none";
    cycloneii_io ix46193z43919 (.padio (o_image1_0_[5]), .datain (nx46193z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix46193z43919.operation_mode = "output";
                 
                 defparam ix46193z43919.output_register_mode = "none";
                 
                 defparam ix46193z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix46193z43919.oe_register_mode = "none";
                 
                 defparam ix46193z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix46193z43919.input_register_mode = "none";
    cycloneii_io ix45196z43919 (.padio (o_image1_0_[4]), .datain (nx45196z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix45196z43919.operation_mode = "output";
                 
                 defparam ix45196z43919.output_register_mode = "none";
                 
                 defparam ix45196z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix45196z43919.oe_register_mode = "none";
                 
                 defparam ix45196z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix45196z43919.input_register_mode = "none";
    cycloneii_io ix44199z43919 (.padio (o_image1_0_[3]), .datain (nx44199z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix44199z43919.operation_mode = "output";
                 
                 defparam ix44199z43919.output_register_mode = "none";
                 
                 defparam ix44199z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix44199z43919.oe_register_mode = "none";
                 
                 defparam ix44199z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix44199z43919.input_register_mode = "none";
    cycloneii_io ix43202z43919 (.padio (o_image1_0_[2]), .datain (nx43202z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix43202z43919.operation_mode = "output";
                 
                 defparam ix43202z43919.output_register_mode = "none";
                 
                 defparam ix43202z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix43202z43919.oe_register_mode = "none";
                 
                 defparam ix43202z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix43202z43919.input_register_mode = "none";
    cycloneii_io ix42205z43919 (.padio (o_image1_0_[1]), .datain (nx42205z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix42205z43919.operation_mode = "output";
                 
                 defparam ix42205z43919.output_register_mode = "none";
                 
                 defparam ix42205z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix42205z43919.oe_register_mode = "none";
                 
                 defparam ix42205z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix42205z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix57374z52923 (.combout (nx57374z1), .dataa (1'b1), .datab (
                         nx57374z2), .datac (mem_q_1_[2]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix57374z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix41208z43919 (.padio (o_image1_0_[0]), .datain (nx41208z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix41208z43919.operation_mode = "output";
                 
                 defparam ix41208z43919.output_register_mode = "none";
                 
                 defparam ix41208z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix41208z43919.oe_register_mode = "none";
                 
                 defparam ix41208z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix41208z43919.input_register_mode = "none";
    cycloneii_io ix43052z43919 (.padio (o_image1_1_[7]), .datain (nx43052z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix43052z43919.operation_mode = "output";
                 
                 defparam ix43052z43919.output_register_mode = "none";
                 
                 defparam ix43052z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix43052z43919.oe_register_mode = "none";
                 
                 defparam ix43052z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix43052z43919.input_register_mode = "none";
    cycloneii_io ix42055z43919 (.padio (o_image1_1_[6]), .datain (nx42055z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix42055z43919.operation_mode = "output";
                 
                 defparam ix42055z43919.output_register_mode = "none";
                 
                 defparam ix42055z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix42055z43919.oe_register_mode = "none";
                 
                 defparam ix42055z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix42055z43919.input_register_mode = "none";
    cycloneii_io ix41058z43919 (.padio (o_image1_1_[5]), .datain (nx41058z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix41058z43919.operation_mode = "output";
                 
                 defparam ix41058z43919.output_register_mode = "none";
                 
                 defparam ix41058z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix41058z43919.oe_register_mode = "none";
                 
                 defparam ix41058z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix41058z43919.input_register_mode = "none";
    cycloneii_io ix40061z43919 (.padio (o_image1_1_[4]), .datain (nx40061z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix40061z43919.operation_mode = "output";
                 
                 defparam ix40061z43919.output_register_mode = "none";
                 
                 defparam ix40061z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix40061z43919.oe_register_mode = "none";
                 
                 defparam ix40061z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix40061z43919.input_register_mode = "none";
    cycloneii_io ix39064z43919 (.padio (o_image1_1_[3]), .datain (nx39064z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix39064z43919.operation_mode = "output";
                 
                 defparam ix39064z43919.output_register_mode = "none";
                 
                 defparam ix39064z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix39064z43919.oe_register_mode = "none";
                 
                 defparam ix39064z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix39064z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix58371z52923 (.combout (nx58371z1), .dataa (1'b1), .datab (
                         nx58371z2), .datac (mem_q_1_[3]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix58371z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix38067z43919 (.padio (o_image1_1_[2]), .datain (nx38067z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix38067z43919.operation_mode = "output";
                 
                 defparam ix38067z43919.output_register_mode = "none";
                 
                 defparam ix38067z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix38067z43919.oe_register_mode = "none";
                 
                 defparam ix38067z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix38067z43919.input_register_mode = "none";
    cycloneii_io ix37070z43919 (.padio (o_image1_1_[1]), .datain (nx37070z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix37070z43919.operation_mode = "output";
                 
                 defparam ix37070z43919.output_register_mode = "none";
                 
                 defparam ix37070z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix37070z43919.oe_register_mode = "none";
                 
                 defparam ix37070z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix37070z43919.input_register_mode = "none";
    cycloneii_io ix36073z43919 (.padio (o_image1_1_[0]), .datain (nx36073z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix36073z43919.operation_mode = "output";
                 
                 defparam ix36073z43919.output_register_mode = "none";
                 
                 defparam ix36073z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix36073z43919.oe_register_mode = "none";
                 
                 defparam ix36073z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix36073z43919.input_register_mode = "none";
    cycloneii_io ix37917z43919 (.padio (o_image1_2_[7]), .datain (nx37917z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix37917z43919.operation_mode = "output";
                 
                 defparam ix37917z43919.output_register_mode = "none";
                 
                 defparam ix37917z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix37917z43919.oe_register_mode = "none";
                 
                 defparam ix37917z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix37917z43919.input_register_mode = "none";
    cycloneii_io ix36920z43919 (.padio (o_image1_2_[6]), .datain (nx36920z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix36920z43919.operation_mode = "output";
                 
                 defparam ix36920z43919.output_register_mode = "none";
                 
                 defparam ix36920z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix36920z43919.oe_register_mode = "none";
                 
                 defparam ix36920z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix36920z43919.input_register_mode = "none";
    cycloneii_io ix35923z43919 (.padio (o_image1_2_[5]), .datain (nx35923z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix35923z43919.operation_mode = "output";
                 
                 defparam ix35923z43919.output_register_mode = "none";
                 
                 defparam ix35923z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix35923z43919.oe_register_mode = "none";
                 
                 defparam ix35923z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix35923z43919.input_register_mode = "none";
    cycloneii_io ix34926z43919 (.padio (o_image1_2_[4]), .datain (nx34926z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix34926z43919.operation_mode = "output";
                 
                 defparam ix34926z43919.output_register_mode = "none";
                 
                 defparam ix34926z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix34926z43919.oe_register_mode = "none";
                 
                 defparam ix34926z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix34926z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix59368z52923 (.combout (nx59368z1), .dataa (1'b1), .datab (
                         nx59368z2), .datac (mem_q_1_[4]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix59368z52923.lut_mask = 16'hf0cc;
    cycloneii_io ix33929z43919 (.padio (o_image1_2_[3]), .datain (nx33929z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix33929z43919.operation_mode = "output";
                 
                 defparam ix33929z43919.output_register_mode = "none";
                 
                 defparam ix33929z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix33929z43919.oe_register_mode = "none";
                 
                 defparam ix33929z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix33929z43919.input_register_mode = "none";
    cycloneii_io ix32932z43919 (.padio (o_image1_2_[2]), .datain (nx32932z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix32932z43919.operation_mode = "output";
                 
                 defparam ix32932z43919.output_register_mode = "none";
                 
                 defparam ix32932z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix32932z43919.oe_register_mode = "none";
                 
                 defparam ix32932z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix32932z43919.input_register_mode = "none";
    cycloneii_io ix31935z43919 (.padio (o_image1_2_[1]), .datain (nx31935z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix31935z43919.operation_mode = "output";
                 
                 defparam ix31935z43919.output_register_mode = "none";
                 
                 defparam ix31935z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix31935z43919.oe_register_mode = "none";
                 
                 defparam ix31935z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix31935z43919.input_register_mode = "none";
    cycloneii_io ix30938z43919 (.padio (o_image1_2_[0]), .datain (nx30938z1), .oe (
                 1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (1'b0), .inclkena (
                 1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam ix30938z43919.operation_mode = "output";
                 
                 defparam ix30938z43919.output_register_mode = "none";
                 
                 defparam ix30938z43919.tie_off_output_clock_enable = "false";
                 
                 defparam ix30938z43919.oe_register_mode = "none";
                 
                 defparam ix30938z43919.tie_off_oe_clock_enable = "false";
                 
                 defparam ix30938z43919.input_register_mode = "none";
    cycloneii_lcell_comb ix60365z52923 (.combout (nx60365z1), .dataa (1'b1), .datab (
                         nx60365z2), .datac (mem_q_1_[5]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix60365z52923.lut_mask = 16'hf0cc;
    cycloneii_lcell_comb ix61362z52923 (.combout (nx61362z1), .dataa (1'b1), .datab (
                         nx61362z2), .datac (mem_q_1_[6]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix61362z52923.lut_mask = 16'hf0cc;
    cycloneii_lcell_comb ix62359z52923 (.combout (nx62359z1), .dataa (1'b1), .datab (
                         nx62359z2), .datac (mem_q_1_[7]), .datad (nx62359z4), .cin (
                         1'b0)) ;
                         defparam ix62359z52923.lut_mask = 16'hf0cc;
    cycloneii_io i_reset_ibuf (.combout (i_reset_int), .padio (i_reset), .datain (
                 1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (
                 1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam i_reset_ibuf.operation_mode = "input";
                 
                 defparam i_reset_ibuf.output_register_mode = "none";
                 
                 defparam i_reset_ibuf.tie_off_output_clock_enable = "false";
                 
                 defparam i_reset_ibuf.oe_register_mode = "none";
                 
                 defparam i_reset_ibuf.tie_off_oe_clock_enable = "false";
                 
                 defparam i_reset_ibuf.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_7_ (.combout (i_pixel_int[7]), .padio (i_pixel[7])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_7_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_7_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_7_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_7_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_7_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_7_.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_6_ (.combout (i_pixel_int[6]), .padio (i_pixel[6])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_6_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_6_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_6_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_6_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_6_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_6_.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_5_ (.combout (i_pixel_int[5]), .padio (i_pixel[5])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_5_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_5_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_5_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_5_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_5_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_5_.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_4_ (.combout (i_pixel_int[4]), .padio (i_pixel[4])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_4_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_4_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_4_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_4_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_4_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_4_.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_3_ (.combout (i_pixel_int[3]), .padio (i_pixel[3])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_3_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_3_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_3_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_3_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_3_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_3_.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_2_ (.combout (i_pixel_int[2]), .padio (i_pixel[2])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_2_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_2_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_2_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_2_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_2_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_2_.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_1_ (.combout (i_pixel_int[1]), .padio (i_pixel[1])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_1_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_1_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_1_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_1_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_1_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_1_.input_register_mode = "none";
    cycloneii_io i_pixel_ibuf_0_ (.combout (i_pixel_int[0]), .padio (i_pixel[0])
                 , .datain (1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1)
                 , .inclk (1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (
                 1'b0)) ;
                 defparam i_pixel_ibuf_0_.operation_mode = "input";
                 
                 defparam i_pixel_ibuf_0_.output_register_mode = "none";
                 
                 defparam i_pixel_ibuf_0_.tie_off_output_clock_enable = "false";
                 defparam i_pixel_ibuf_0_.oe_register_mode = "none";
                 
                 defparam i_pixel_ibuf_0_.tie_off_oe_clock_enable = "false";
                 defparam i_pixel_ibuf_0_.input_register_mode = "none";
    cycloneii_io i_clock_ibuf (.combout (i_clock_int), .padio (i_clock), .datain (
                 1'b0), .oe (1'b1), .outclk (1'b0), .outclkena (1'b1), .inclk (
                 1'b0), .inclkena (1'b1), .areset (1'b0), .sreset (1'b0)) ;
                 
                 defparam i_clock_ibuf.operation_mode = "input";
                 
                 defparam i_clock_ibuf.output_register_mode = "none";
                 
                 defparam i_clock_ibuf.tie_off_output_clock_enable = "false";
                 
                 defparam i_clock_ibuf.oe_register_mode = "none";
                 
                 defparam i_clock_ibuf.tie_off_oe_clock_enable = "false";
                 
                 defparam i_clock_ibuf.input_register_mode = "none";
    cycloneii_lcell_comb ix8852z52927 (.combout (nx8852z5), .dataa (column[3]), 
                         .datab (column[2]), .datac (1'b1), .datad (1'b1), .cin (
                         1'b0)) ;
                         defparam ix8852z52927.lut_mask = 16'h8888;
    cycloneii_lcell_comb ix41103z52924 (.combout (nx41103z2), .dataa (
                         mem_wrn_current[2]), .datab (mem_wrn_current[1]), .datac (
                         mem_wrn_current[0]), .datad (i_valid_int), .cin (1'b0)
                         ) ;
                         defparam ix41103z52924.lut_mask = 16'h01ff;
    cycloneii_lcell_comb ix41103z52925 (.combout (nx41103z3), .dataa (
                         first_bubble), .datab (nx8852z3), .datac (i_valid_int)
                         , .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix41103z52925.lut_mask = 16'h0707;
    cycloneii_lcell_comb ix60567z52928 (.combout (nx60567z6), .dataa (column[3])
                         , .datab (column[2]), .datac (column[1]), .datad (1'b1)
                         , .cin (1'b0)) ;
                         
                         defparam ix60567z52928.lut_mask = 16'hfefe;
    cycloneii_lcell_comb ix62359z52925 (.combout (nx62359z3), .dataa (
                         mem_wrn_current[1]), .datab (mem_wrn_current[0]), .datac (
                         nx60567z2), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix62359z52925.lut_mask = 16'hd5d5;
    cycloneii_lcell_comb ix63578z52926 (.combout (nx63578z3), .dataa (
                         mem_wrn_current[1]), .datab (mem_wrn_current[0]), .datac (
                         nx60567z2), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix63578z52926.lut_mask = 16'hb3b3;
    cycloneii_lcell_comb ix60567z52927 (.combout (nx60567z5), .dataa (column[6])
                         , .datab (column[5]), .datac (column[4]), .datad (
                         nx60567z2), .cin (1'b0)) ;
                         
                         defparam ix60567z52927.lut_mask = 16'hfe00;
    cycloneii_lcell_comb ix60567z52926 (.combout (nx60567z4), .dataa (
                         o_valid_dup0), .datab (column[7]), .datac (nx60567z2), 
                         .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix60567z52926.lut_mask = 16'heaea;
    cycloneii_lcell_comb ix60567z52925 (.combout (nx60567z3), .dataa (row[4]), .datab (
                         row[3]), .datac (row[2]), .datad (row[1]), .cin (1'b0)
                         ) ;
                         defparam ix60567z52925.lut_mask = 16'hfffe;
    cycloneii_lcell_comb ix8852z52929 (.combout (nx8852z7), .dataa (row[3]), .datab (
                         row[2]), .datac (row[1]), .datad (row[0]), .cin (1'b0)
                         ) ;
                         defparam ix8852z52929.lut_mask = 16'h8000;
    cycloneii_lcell_comb ix8852z52928 (.combout (nx8852z6), .dataa (row[7]), .datab (
                         row[6]), .datac (row[5]), .datad (row[4]), .cin (1'b0)
                         ) ;
                         defparam ix8852z52928.lut_mask = 16'h8000;
    cycloneii_lcell_comb ix8852z52926 (.combout (nx8852z4), .dataa (column[7]), 
                         .datab (column[6]), .datac (column[5]), .datad (
                         column[4]), .cin (1'b0)) ;
                         
                         defparam ix8852z52926.lut_mask = 16'h8000;
    cycloneii_lcell_comb ix39109z52924 (.combout (nx39109z2), .dataa (nx8852z2)
                         , .datab (i_reset_int), .datac (nx41103z3), .datad (
                         nx41103z2), .cin (1'b0)) ;
                         
                         defparam ix39109z52924.lut_mask = 16'hefee;
    cycloneii_lcell_comb ix62359z52924 (.combout (nx62359z2), .dataa (
                         buffer2_4n2ss1[7]), .datab (mem_q_2_[7]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix62359z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix61362z52924 (.combout (nx61362z2), .dataa (
                         buffer2_4n2ss1[6]), .datab (mem_q_2_[6]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix61362z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix60365z52924 (.combout (nx60365z2), .dataa (
                         buffer2_4n2ss1[5]), .datab (mem_q_2_[5]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix60365z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix59368z52924 (.combout (nx59368z2), .dataa (
                         buffer2_4n2ss1[4]), .datab (mem_q_2_[4]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix59368z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix58371z52924 (.combout (nx58371z2), .dataa (
                         buffer2_4n2ss1[3]), .datab (mem_q_2_[3]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix58371z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix57374z52924 (.combout (nx57374z2), .dataa (
                         buffer2_4n2ss1[2]), .datab (mem_q_2_[2]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix57374z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix56377z52924 (.combout (nx56377z2), .dataa (
                         buffer2_4n2ss1[1]), .datab (mem_q_2_[1]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix56377z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix55380z52924 (.combout (nx55380z2), .dataa (
                         buffer2_4n2ss1[0]), .datab (mem_q_2_[0]), .datac (
                         nx62359z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix55380z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix63578z52924 (.combout (nx63578z2), .dataa (
                         buffer2_4n2ss1[7]), .datab (mem_q_2_[7]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix63578z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix64575z52924 (.combout (nx64575z2), .dataa (
                         buffer2_4n2ss1[6]), .datab (mem_q_2_[6]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix64575z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix36z52924 (.combout (nx36z2), .dataa (
                         buffer2_4n2ss1[5]), .datab (mem_q_2_[5]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix36z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix1033z52924 (.combout (nx1033z2), .dataa (
                         buffer2_4n2ss1[4]), .datab (mem_q_2_[4]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix1033z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix2030z52924 (.combout (nx2030z2), .dataa (
                         buffer2_4n2ss1[3]), .datab (mem_q_2_[3]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix2030z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix3027z52924 (.combout (nx3027z2), .dataa (
                         buffer2_4n2ss1[2]), .datab (mem_q_2_[2]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix3027z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix4024z52924 (.combout (nx4024z2), .dataa (
                         buffer2_4n2ss1[1]), .datab (mem_q_2_[1]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix4024z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix5021z52924 (.combout (nx5021z2), .dataa (
                         buffer2_4n2ss1[0]), .datab (mem_q_2_[0]), .datac (
                         nx63578z3), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix5021z52924.lut_mask = 16'hcaca;
    cycloneii_lcell_comb ix60567z52923 (.combout (nx60567z1), .dataa (nx60567z2)
                         , .datab (nx60567z4), .datac (nx60567z5), .datad (
                         nx60567z6), .cin (1'b0)) ;
                         
                         defparam ix60567z52923.lut_mask = 16'hfefc;
    cycloneii_lcell_comb ix8852z52925 (.combout (nx8852z3), .dataa (column[1]), 
                         .datab (column[0]), .datac (nx8852z4), .datad (nx8852z5
                         ), .cin (1'b0)) ;
                         
                         defparam ix8852z52925.lut_mask = 16'h8000;
    cycloneii_lcell_comb ix62359z52926 (.combout (nx62359z4), .dataa (
                         mem_wrn_current[1]), .datab (mem_wrn_current[0]), .datac (
                         nx60567z2), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix62359z52926.lut_mask = 16'h1515;
    cycloneii_lcell_comb ix63578z52927 (.combout (nx63578z4), .dataa (
                         mem_wrn_current[1]), .datab (mem_wrn_current[0]), .datac (
                         nx60567z2), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix63578z52927.lut_mask = 16'h1313;
    cycloneii_lcell_comb ix41103z52926 (.combout (nx41103z4), .dataa (nx8852z1)
                         , .datab (i_valid_int), .datac (nx41103z3), .datad (
                         nx41103z2), .cin (1'b0)) ;
                         
                         defparam ix41103z52926.lut_mask = 16'haeaa;
    cycloneii_lcell_comb ix33254z52923 (.combout (nx33254z1), .dataa (busySignal
                         ), .datab (i_valid_int), .datac (1'b1), .datad (1'b1), 
                         .cin (1'b0)) ;
                         
                         defparam ix33254z52923.lut_mask = 16'heeee;
    cycloneii_lcell_comb ix8852z52924 (.combout (nx8852z2), .dataa (first_bubble
                         ), .datab (nx8852z3), .datac (nx8852z6), .datad (
                         nx8852z7), .cin (1'b0)) ;
                         
                         defparam ix8852z52924.lut_mask = 16'h8000;
    cycloneii_lcell_comb ix60567z52924 (.combout (nx60567z2), .dataa (row[7]), .datab (
                         row[6]), .datac (row[5]), .datad (nx60567z3), .cin (
                         1'b0)) ;
                         defparam ix60567z52924.lut_mask = 16'hfffe;
    cycloneii_lcell_comb ix5021z52925 (.combout (buffer2_4n2ss1[0]), .dataa (
                         nx60567z2), .datab (mem_q_1_[0]), .datac (
                         i_pixel_int[0]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix5021z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix4024z52925 (.combout (buffer2_4n2ss1[1]), .dataa (
                         nx60567z2), .datab (mem_q_1_[1]), .datac (
                         i_pixel_int[1]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix4024z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix3027z52925 (.combout (buffer2_4n2ss1[2]), .dataa (
                         nx60567z2), .datab (mem_q_1_[2]), .datac (
                         i_pixel_int[2]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix3027z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix2030z52925 (.combout (buffer2_4n2ss1[3]), .dataa (
                         nx60567z2), .datab (mem_q_1_[3]), .datac (
                         i_pixel_int[3]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix2030z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix1033z52925 (.combout (buffer2_4n2ss1[4]), .dataa (
                         nx60567z2), .datab (mem_q_1_[4]), .datac (
                         i_pixel_int[4]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix1033z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix36z52925 (.combout (buffer2_4n2ss1[5]), .dataa (
                         nx60567z2), .datab (mem_q_1_[5]), .datac (
                         i_pixel_int[5]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix36z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix64575z52925 (.combout (buffer2_4n2ss1[6]), .dataa (
                         nx60567z2), .datab (mem_q_1_[6]), .datac (
                         i_pixel_int[6]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix64575z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix63578z52925 (.combout (buffer2_4n2ss1[7]), .dataa (
                         nx60567z2), .datab (mem_q_1_[7]), .datac (
                         i_pixel_int[7]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix63578z52925.lut_mask = 16'hd8d8;
    cycloneii_lcell_comb ix15763z52925 (.combout (nx15763z3), .dataa (nx15763z4)
                         , .datab (nx8852z2), .datac (i_valid_int), .datad (
                         i_reset_int), .cin (1'b0)) ;
                         
                         defparam ix15763z52925.lut_mask = 16'h0010;
    cycloneii_lcell_comb ix8852z52930 (.combout (not_rtlc3_X_0_n252), .dataa (
                         first_bubble), .datab (nx8852z3), .datac (i_valid_int)
                         , .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix8852z52930.lut_mask = 16'h0808;
    cycloneii_lcell_comb ix15763z52926 (.combout (nx15763z4), .dataa (
                         mem_wrn_current[2]), .datab (mem_wrn_current[1]), .datac (
                         mem_wrn_current[0]), .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix15763z52926.lut_mask = 16'hfefe;
    cycloneii_lcell_comb ix8852z52923 (.combout (nx8852z1), .dataa (nx8852z2), .datab (
                         i_reset_int), .datac (1'b1), .datad (1'b1), .cin (1'b0)
                         ) ;
                         defparam ix8852z52923.lut_mask = 16'heeee;
    cycloneii_lcell_comb ix47893z52923 (.combout (o_mode_dup0[0]), .dataa (
                         busySignal), .datab (busySignalDelayed), .datac (
                         i_valid_int), .datad (i_reset_int), .cin (1'b0)) ;
                         
                         defparam ix47893z52923.lut_mask = 16'hfffe;
    cycloneii_lcell_comb ix50245z52923 (.combout (nx50245z1), .dataa (
                         i_pixel_int[0]), .datab (mem_q_2_[0]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix50245z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix51242z52923 (.combout (nx51242z1), .dataa (
                         i_pixel_int[1]), .datab (mem_q_2_[1]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix51242z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix52239z52923 (.combout (nx52239z1), .dataa (
                         i_pixel_int[2]), .datab (mem_q_2_[2]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix52239z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix53236z52923 (.combout (nx53236z1), .dataa (
                         i_pixel_int[3]), .datab (mem_q_2_[3]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix53236z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix54233z52923 (.combout (nx54233z1), .dataa (
                         i_pixel_int[4]), .datab (mem_q_2_[4]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix54233z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix55230z52923 (.combout (nx55230z1), .dataa (
                         i_pixel_int[5]), .datab (mem_q_2_[5]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix55230z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix56227z52923 (.combout (nx56227z1), .dataa (
                         i_pixel_int[6]), .datab (mem_q_2_[6]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix56227z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix57224z52923 (.combout (nx57224z1), .dataa (
                         i_pixel_int[7]), .datab (mem_q_2_[7]), .datac (
                         nx60567z2), .datad (mem_wrn_current[2]), .cin (1'b0)) ;
                         
                         defparam ix57224z52923.lut_mask = 16'haaac;
    cycloneii_lcell_comb ix39109z52925 (.combout (nx39109z3), .dataa (
                         i_valid_int), .datab (mem_wrn_current[0]), .datac (
                         mem_wrn_current[1]), .datad (mem_wrn_current[2]), .cin (
                         1'b0)) ;
                         defparam ix39109z52925.lut_mask = 16'h0002;
    cycloneii_lcell_comb ix41103z52923 (.combout (nx41103z1), .dataa (nx41103z2)
                         , .datab (nx41103z3), .datac (i_reset_int), .datad (
                         nx8852z2), .cin (1'b0)) ;
                         
                         defparam ix41103z52923.lut_mask = 16'hfff2;
    cycloneii_lcell_comb ix16760z52923 (.combout (nx16760z1), .dataa (nx41103z2)
                         , .datab (i_reset_int), .datac (nx8852z2), .datad (1'b1
                         ), .cin (1'b0)) ;
                         
                         defparam ix16760z52923.lut_mask = 16'hfefe;
    cycloneii_lcell_comb ix15763z52924 (.combout (nx15763z2), .dataa (
                         i_valid_int), .datab (i_reset_int), .datac (nx8852z2), 
                         .datad (1'b1), .cin (1'b0)) ;
                         
                         defparam ix15763z52924.lut_mask = 16'hfdfd;
    cycloneii_lcell_comb ix47386z52923 (.combout (nx47386z1), .dataa (nx8852z3)
                         , .datab (first_bubble), .datac (i_reset_int), .datad (
                         nx8852z2), .cin (1'b0)) ;
                         
                         defparam ix47386z52923.lut_mask = 16'hfff8;
endmodule


module ram_dq_8_2 ( wr_data1, rd_data1, addr1, wr_clk1, rd_clk1, wr_ena1, 
                    rd_ena1, ena1, rst1, regce1 ) ;

    input [7:0]wr_data1 ;
    output [7:0]rd_data1 ;
    input [7:0]addr1 ;
    input wr_clk1 ;
    input rd_clk1 ;
    input wr_ena1 ;
    input rd_ena1 ;
    input ena1 ;
    input rst1 ;
    input regce1 ;

    wire ena1_rename637;



    altsyncram ix64056z29483 (.data_a ({wr_data1[7],wr_data1[6],wr_data1[5],
               wr_data1[4],wr_data1[3],wr_data1[2],wr_data1[1],wr_data1[0]}), .address_a (
               {addr1[7],addr1[6],addr1[5],addr1[4],addr1[3],addr1[2],addr1[1],
               addr1[0]}), .wren_a (wr_ena1), .clock0 (wr_clk1), .clocken0 (
               ena1_rename637), .q_a ({rd_data1[7],rd_data1[6],rd_data1[5],
               rd_data1[4],rd_data1[3],rd_data1[2],rd_data1[1],rd_data1[0]})) ;
               
               defparam ix64056z29483.width_a = 8;
               
               defparam ix64056z29483.widthad_a = 8;
               
               defparam ix64056z29483.numwords_a = 256;
               
               defparam ix64056z29483.outdata_reg_a = "UNREGISTERED";
               
               defparam ix64056z29483.address_aclr_a = "NONE";
               
               defparam ix64056z29483.outdata_aclr_a = "NONE";
               
               defparam ix64056z29483.indata_aclr_a = "NONE";
               
               defparam ix64056z29483.wrcontrol_aclr_a = "NONE";
               
               defparam ix64056z29483.byteena_aclr_a = "NONE";
               
               defparam ix64056z29483.width_byteena_a = 1;
               
               defparam ix64056z29483.width_b = 8;
               
               defparam ix64056z29483.widthad_b = 8;
               
               defparam ix64056z29483.numwords_b = 256;
               
               defparam ix64056z29483.rdcontrol_reg_b = "CLOCK1";
               
               defparam ix64056z29483.address_reg_b = "CLOCK1";
               
               defparam ix64056z29483.outdata_reg_b = "UNREGISTERED";
               
               defparam ix64056z29483.outdata_aclr_b = "NONE";
               
               defparam ix64056z29483.rdcontrol_aclr_b = "NONE";
               
               defparam ix64056z29483.indata_reg_b = "CLOCK1";
               
               defparam ix64056z29483.wrcontrol_wraddress_reg_b = "CLOCK1";
               
               defparam ix64056z29483.byteena_reg_b = "CLOCK1";
               
               defparam ix64056z29483.indata_aclr_b = "NONE";
               
               defparam ix64056z29483.wrcontrol_aclr_b = "NONE";
               
               defparam ix64056z29483.byteena_aclr_b = "NONE";
               
               defparam ix64056z29483.width_byteena_b = 1;
               
               defparam ix64056z29483.address_aclr_b = "NONE";
               
               defparam ix64056z29483.operation_mode = "SINGLE_PORT";
               
               defparam ix64056z29483.byte_size = 8;
               
               defparam ix64056z29483.read_during_write_mode_mixed_ports = "DONT_CARE";
               
               defparam ix64056z29483.ram_block_type = "AUTO";
               
               defparam ix64056z29483.init_file = "UNUSED";
               
               defparam ix64056z29483.init_file_layout = "UNUSED";
               
               defparam ix64056z29483.maximum_depth = 0;
               
               defparam ix64056z29483.intended_device_family = "Stratix";
               
               defparam ix64056z29483.lpm_hint = "UNUSED";
               
               defparam ix64056z29483.lpm_type = "altsyncram";
    assign ena1_rename637 = 1 ;
endmodule


module ram_dq_8_1 ( wr_data1, rd_data1, addr1, wr_clk1, rd_clk1, wr_ena1, 
                    rd_ena1, ena1, rst1, regce1 ) ;

    input [7:0]wr_data1 ;
    output [7:0]rd_data1 ;
    input [7:0]addr1 ;
    input wr_clk1 ;
    input rd_clk1 ;
    input wr_ena1 ;
    input rd_ena1 ;
    input ena1 ;
    input rst1 ;
    input regce1 ;

    wire ena1_rename607;



    altsyncram ix64056z29482 (.data_a ({wr_data1[7],wr_data1[6],wr_data1[5],
               wr_data1[4],wr_data1[3],wr_data1[2],wr_data1[1],wr_data1[0]}), .address_a (
               {addr1[7],addr1[6],addr1[5],addr1[4],addr1[3],addr1[2],addr1[1],
               addr1[0]}), .wren_a (wr_ena1), .clock0 (wr_clk1), .clocken0 (
               ena1_rename607), .q_a ({rd_data1[7],rd_data1[6],rd_data1[5],
               rd_data1[4],rd_data1[3],rd_data1[2],rd_data1[1],rd_data1[0]})) ;
               
               defparam ix64056z29482.width_a = 8;
               
               defparam ix64056z29482.widthad_a = 8;
               
               defparam ix64056z29482.numwords_a = 256;
               
               defparam ix64056z29482.outdata_reg_a = "UNREGISTERED";
               
               defparam ix64056z29482.address_aclr_a = "NONE";
               
               defparam ix64056z29482.outdata_aclr_a = "NONE";
               
               defparam ix64056z29482.indata_aclr_a = "NONE";
               
               defparam ix64056z29482.wrcontrol_aclr_a = "NONE";
               
               defparam ix64056z29482.byteena_aclr_a = "NONE";
               
               defparam ix64056z29482.width_byteena_a = 1;
               
               defparam ix64056z29482.width_b = 8;
               
               defparam ix64056z29482.widthad_b = 8;
               
               defparam ix64056z29482.numwords_b = 256;
               
               defparam ix64056z29482.rdcontrol_reg_b = "CLOCK1";
               
               defparam ix64056z29482.address_reg_b = "CLOCK1";
               
               defparam ix64056z29482.outdata_reg_b = "UNREGISTERED";
               
               defparam ix64056z29482.outdata_aclr_b = "NONE";
               
               defparam ix64056z29482.rdcontrol_aclr_b = "NONE";
               
               defparam ix64056z29482.indata_reg_b = "CLOCK1";
               
               defparam ix64056z29482.wrcontrol_wraddress_reg_b = "CLOCK1";
               
               defparam ix64056z29482.byteena_reg_b = "CLOCK1";
               
               defparam ix64056z29482.indata_aclr_b = "NONE";
               
               defparam ix64056z29482.wrcontrol_aclr_b = "NONE";
               
               defparam ix64056z29482.byteena_aclr_b = "NONE";
               
               defparam ix64056z29482.width_byteena_b = 1;
               
               defparam ix64056z29482.address_aclr_b = "NONE";
               
               defparam ix64056z29482.operation_mode = "SINGLE_PORT";
               
               defparam ix64056z29482.byte_size = 8;
               
               defparam ix64056z29482.read_during_write_mode_mixed_ports = "DONT_CARE";
               
               defparam ix64056z29482.ram_block_type = "AUTO";
               
               defparam ix64056z29482.init_file = "UNUSED";
               
               defparam ix64056z29482.init_file_layout = "UNUSED";
               
               defparam ix64056z29482.maximum_depth = 0;
               
               defparam ix64056z29482.intended_device_family = "Stratix";
               
               defparam ix64056z29482.lpm_hint = "UNUSED";
               
               defparam ix64056z29482.lpm_type = "altsyncram";
    assign ena1_rename607 = 1 ;
endmodule


module ram_dq_8_0 ( wr_data1, rd_data1, addr1, wr_clk1, rd_clk1, wr_ena1, 
                    rd_ena1, ena1, rst1, regce1 ) ;

    input [7:0]wr_data1 ;
    output [7:0]rd_data1 ;
    input [7:0]addr1 ;
    input wr_clk1 ;
    input rd_clk1 ;
    input wr_ena1 ;
    input rd_ena1 ;
    input ena1 ;
    input rst1 ;
    input regce1 ;

    wire ena1_rename577;



    altsyncram ix64056z29481 (.data_a ({wr_data1[7],wr_data1[6],wr_data1[5],
               wr_data1[4],wr_data1[3],wr_data1[2],wr_data1[1],wr_data1[0]}), .address_a (
               {addr1[7],addr1[6],addr1[5],addr1[4],addr1[3],addr1[2],addr1[1],
               addr1[0]}), .wren_a (wr_ena1), .clock0 (wr_clk1), .clocken0 (
               ena1_rename577), .q_a ({rd_data1[7],rd_data1[6],rd_data1[5],
               rd_data1[4],rd_data1[3],rd_data1[2],rd_data1[1],rd_data1[0]})) ;
               
               defparam ix64056z29481.width_a = 8;
               
               defparam ix64056z29481.widthad_a = 8;
               
               defparam ix64056z29481.numwords_a = 256;
               
               defparam ix64056z29481.outdata_reg_a = "UNREGISTERED";
               
               defparam ix64056z29481.address_aclr_a = "NONE";
               
               defparam ix64056z29481.outdata_aclr_a = "NONE";
               
               defparam ix64056z29481.indata_aclr_a = "NONE";
               
               defparam ix64056z29481.wrcontrol_aclr_a = "NONE";
               
               defparam ix64056z29481.byteena_aclr_a = "NONE";
               
               defparam ix64056z29481.width_byteena_a = 1;
               
               defparam ix64056z29481.width_b = 8;
               
               defparam ix64056z29481.widthad_b = 8;
               
               defparam ix64056z29481.numwords_b = 256;
               
               defparam ix64056z29481.rdcontrol_reg_b = "CLOCK1";
               
               defparam ix64056z29481.address_reg_b = "CLOCK1";
               
               defparam ix64056z29481.outdata_reg_b = "UNREGISTERED";
               
               defparam ix64056z29481.outdata_aclr_b = "NONE";
               
               defparam ix64056z29481.rdcontrol_aclr_b = "NONE";
               
               defparam ix64056z29481.indata_reg_b = "CLOCK1";
               
               defparam ix64056z29481.wrcontrol_wraddress_reg_b = "CLOCK1";
               
               defparam ix64056z29481.byteena_reg_b = "CLOCK1";
               
               defparam ix64056z29481.indata_aclr_b = "NONE";
               
               defparam ix64056z29481.wrcontrol_aclr_b = "NONE";
               
               defparam ix64056z29481.byteena_aclr_b = "NONE";
               
               defparam ix64056z29481.width_byteena_b = 1;
               
               defparam ix64056z29481.address_aclr_b = "NONE";
               
               defparam ix64056z29481.operation_mode = "SINGLE_PORT";
               
               defparam ix64056z29481.byte_size = 8;
               
               defparam ix64056z29481.read_during_write_mode_mixed_ports = "DONT_CARE";
               
               defparam ix64056z29481.ram_block_type = "AUTO";
               
               defparam ix64056z29481.init_file = "UNUSED";
               
               defparam ix64056z29481.init_file_layout = "UNUSED";
               
               defparam ix64056z29481.maximum_depth = 0;
               
               defparam ix64056z29481.intended_device_family = "Stratix";
               
               defparam ix64056z29481.lpm_hint = "UNUSED";
               
               defparam ix64056z29481.lpm_type = "altsyncram";
    assign ena1_rename577 = 1 ;
endmodule


module modgen_counter_8_1 ( clock, q, clk_en, aclear, sload, data, aset, sclear, 
                            updn, cnt_en, p_rtlc3n121, p_i_valid_int ) ;

    input clock ;
    output [7:0]q ;
    input clk_en ;
    input aclear ;
    input sload ;
    input [7:0]data ;
    input aset ;
    input sclear ;
    input updn ;
    input cnt_en ;
    input p_rtlc3n121 ;
    input p_i_valid_int ;

    wire nx57253z3, nx51271z1, nx58250z14, nx52268z1, nx58250z12, nx53265z1, 
         nx58250z10, nx54262z1, nx58250z8, nx55259z1, nx58250z6, nx56256z1, 
         nx58250z4, nx57253z1, nx58250z2, nx58250z1, 
         nx_modgen_counter_8_1_vcc_net;
    wire [43:0] xmplr_dummy ;




    cycloneii_lcell_ff reg_q_7_ (.regout (q[7]), .datain (nx58250z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_6_ (.regout (q[6]), .datain (nx57253z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_5_ (.regout (q[5]), .datain (nx56256z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_4_ (.regout (q[4]), .datain (nx55259z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_3_ (.regout (q[3]), .datain (nx54262z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_2_ (.regout (q[2]), .datain (nx53265z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_1_ (.regout (q[1]), .datain (nx52268z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_0_ (.regout (q[0]), .datain (nx51271z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_comb ix58250z52929 (.combout (nx53265z1), .cout (nx58250z10)
                         , .dataa (q[2]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (nx58250z12)) ;
                         
                         defparam ix58250z52929.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52929.sum_lutc_input = "cin";
    assign nx_modgen_counter_8_1_vcc_net = 1 ;
    cycloneii_lcell_comb ix58250z52923 (.combout (nx58250z1), .dataa (q[7]), .datab (
                         1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (nx58250z2)) ;
                         
                         defparam ix58250z52923.lut_mask = 16'h5a00;
                         
                         defparam ix58250z52923.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52925 (.combout (nx57253z1), .cout (nx58250z2)
                         , .dataa (q[6]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (nx58250z4)) ;
                         
                         defparam ix58250z52925.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52925.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52930 (.combout (nx52268z1), .cout (nx58250z12)
                         , .dataa (q[1]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (nx58250z14)) ;
                         
                         defparam ix58250z52930.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52930.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52926 (.combout (nx56256z1), .cout (nx58250z4)
                         , .dataa (q[5]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (nx58250z6)) ;
                         
                         defparam ix58250z52926.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52926.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52927 (.combout (nx55259z1), .cout (nx58250z6)
                         , .dataa (q[4]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (nx58250z8)) ;
                         
                         defparam ix58250z52927.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52927.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52928 (.combout (nx54262z1), .cout (nx58250z8)
                         , .dataa (q[3]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (nx58250z10)) ;
                         
                         defparam ix58250z52928.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52928.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52931 (.combout (nx51271z1), .cout (nx58250z14)
                         , .dataa (q[0]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_1_vcc_net), .cin (1'b0)) ;
                         
                         defparam ix58250z52931.lut_mask = 16'h55aa;
    cycloneii_lcell_comb ix57253z52923 (.combout (nx57253z3), .dataa (cnt_en), .datab (
                         sclear), .datac (p_i_valid_int), .datad (p_rtlc3n121), 
                         .cin (1'b0)) ;
                         
                         defparam ix57253z52923.lut_mask = 16'hee0e;
endmodule


module modgen_counter_8_0 ( clock, q, clk_en, aclear, sload, data, aset, sclear, 
                            updn, cnt_en, p_rtlc6n55, p_i_reset_int ) ;

    input clock ;
    output [7:0]q ;
    input clk_en ;
    input aclear ;
    input sload ;
    input [7:0]data ;
    input aset ;
    input sclear ;
    input updn ;
    input cnt_en ;
    input p_rtlc6n55 ;
    input p_i_reset_int ;

    wire nx57253z3, nx51271z1, nx58250z14, nx52268z1, nx58250z12, nx53265z1, 
         nx58250z10, nx54262z1, nx58250z8, nx55259z1, nx58250z6, nx56256z1, 
         nx58250z4, nx57253z1, nx58250z2, nx58250z1, 
         nx_modgen_counter_8_0_vcc_net;
    wire [44:0] xmplr_dummy ;




    cycloneii_lcell_ff reg_q_7_ (.regout (q[7]), .datain (nx58250z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_6_ (.regout (q[6]), .datain (nx57253z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_5_ (.regout (q[5]), .datain (nx56256z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_4_ (.regout (q[4]), .datain (nx55259z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_3_ (.regout (q[3]), .datain (nx54262z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_2_ (.regout (q[2]), .datain (nx53265z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_1_ (.regout (q[1]), .datain (nx52268z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_ff reg_q_0_ (.regout (q[0]), .datain (nx51271z1), .sdata (
                       1'b0), .clk (clock), .ena (nx57253z3), .aclr (1'b0), .sclr (
                       sclear), .sload (1'b0)) ;
    cycloneii_lcell_comb ix58250z52929 (.combout (nx53265z1), .cout (nx58250z10)
                         , .dataa (q[2]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (nx58250z12)) ;
                         
                         defparam ix58250z52929.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52929.sum_lutc_input = "cin";
    assign nx_modgen_counter_8_0_vcc_net = 1 ;
    cycloneii_lcell_comb ix58250z52923 (.combout (nx58250z1), .dataa (q[7]), .datab (
                         1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (nx58250z2)) ;
                         
                         defparam ix58250z52923.lut_mask = 16'h5a00;
                         
                         defparam ix58250z52923.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52925 (.combout (nx57253z1), .cout (nx58250z2)
                         , .dataa (q[6]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (nx58250z4)) ;
                         
                         defparam ix58250z52925.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52925.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52930 (.combout (nx52268z1), .cout (nx58250z12)
                         , .dataa (q[1]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (nx58250z14)) ;
                         
                         defparam ix58250z52930.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52930.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52926 (.combout (nx56256z1), .cout (nx58250z4)
                         , .dataa (q[5]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (nx58250z6)) ;
                         
                         defparam ix58250z52926.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52926.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52927 (.combout (nx55259z1), .cout (nx58250z6)
                         , .dataa (q[4]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (nx58250z8)) ;
                         
                         defparam ix58250z52927.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52927.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52928 (.combout (nx54262z1), .cout (nx58250z8)
                         , .dataa (q[3]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (nx58250z10)) ;
                         
                         defparam ix58250z52928.lut_mask = 16'h5aa0;
                         
                         defparam ix58250z52928.sum_lutc_input = "cin";
    cycloneii_lcell_comb ix58250z52931 (.combout (nx51271z1), .cout (nx58250z14)
                         , .dataa (q[0]), .datab (1'b1), .datac (1'b1), .datad (
                         nx_modgen_counter_8_0_vcc_net), .cin (1'b0)) ;
                         
                         defparam ix58250z52931.lut_mask = 16'h55aa;
    cycloneii_lcell_comb ix57253z52923 (.combout (nx57253z3), .dataa (cnt_en), .datab (
                         p_i_reset_int), .datac (p_rtlc6n55), .datad (1'b1), .cin (
                         1'b0)) ;
                         defparam ix57253z52923.lut_mask = 16'hfefe;
endmodule

